//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
lX0avB35pFh9RnwDi20I6/Zqm0iWbH4P47tWqxdP+FtA9fGQZ116cq0UjQ3Fig33
MMtZbBG5oG6ZPUrVrkRMF23L/geB0VmFyL7Dac/vOU13WR1K+tWi8pOnDE8JABmS
1NizoNHr8pNd6wLaAqhG/ccm6gyuJyscN1eIu1YN3UxEFfXvi547fXHchNn21mbr
ZGcp17qX/a0q98S8TBrrdZH2y28ErxDdgrLjRsRzQ9zFqE2lfrfiuGz+3rkVpjA3
Qixljiz04VUzDIzU/uN+0nTqp9pHPqjATmIgIRomiq0tJHHXXpxpqjwTi2ZgK/7/
6mC4fReLeP7Xz9LCJYDK8g==
//pragma protect end_key_block
//pragma protect digest_block
hAhA0xBsRYo4Hl1OZKi25fo0AZI=
//pragma protect end_digest_block
//pragma protect data_block
DUOYrF/w6oL3B3TdCT6FB1mhZEgs0KA6j5qO/OkJA6vZkcC6ScprO6py/QCK/hk1
sD4BVxscP+yVWe9ippORqzK97k0ZK5hma9XNwzQ/pebtEfr6krEBddPYRtp3cV+C
O86o+Xho33rMiOxbiBScCPn9GIVgKKse6I0livLpaP3SiIKkMHvBi19MAWS9DsPv
2lsJk1Eaq+IPHzSRAQ1L6w90SJ/k9Ff4PeyKgLHfNpNLqQg0K6RKUTnjUUbqgApQ
HC7rD7dmQwz/TMRO6SlB5/Cm3gc+tyaY0kb6XEyJYLZNzHhqf2gPb+7i+2DG3bH/
RrdrtJeeoRaOHeq87fM9w+mZ+PRS42M0D7MdFADN6KS0fb0LKt5sDaE9swL8ssmS
nlpRHao7JpboIdlL8slgQcVFuTD0JWH5ppQCxYQPk1t4G69oYnPERtBUpZ/RWUbP
gmKFG+NGM6eUS+9wh04RZFyROGMSRXN1yGOGZ3dXQv7jAlm+aHUOJXdTMs6gDbHh
oRt+geZEf7HPr7ipivSakDC+dhC+h2p/izlpTyOurpZrIp+Fka+efH+HjQ3k7qNL
AiyyliHaUxGQ/dvylqyNz+w/drOMOcSUIH0uHthbH6+K7RQ9mNe0snX98PEAEw0v
tklxzf63bIgGPHhPwL5S2FZ10LPmkZujBlj5fSd/ipZ9AcBZBKwsgvvKR3FUkzCb
XA6GKi0EjTVey39hpQqtVw2W1do3yslhmxk3+eR3a8ShXemBUzyueztcHqi1sSyy
+nxe8hUl/IUV6G23D42wpJhRfEKgzueXmoYMLQ0ID+fJqz2Jr1mi+jnSMx4myhL2
No2Oi/B2qVxB2ZL8T0QJnUmES7Q3QXmaxgqcON/baheMjY914Rb6HkdCdbRHWGLH
B6RsWleEkob8bZL1qOEYXWUUYsWsvdZ94SoHV4THC0xP2t+P8crDfsUyluV4Fk2S
g7KaRwCXbEmyzQysucTl2gjLAXaIefPzQMsod3tq2zfpChNxPvm5kfubVAfL9D83
BVZR9a+ZshxJbck7JH70jzuO0XK/bbBG4hbpI0UVdAJNjLD2Sk5+n9iCIpEdGP6v
OBilEMlxUmTB6uY+5ti06gOudgd9W0KZ7ueBlU4dOI3NWTSA3xZf5AJShj5Oio6w
80dVUrmZjoawnMcsSmzpXbbNSAd8MJ454yEZr2dABJjjP8XVUCsLkRlnwWJj5lQl
XSk78aahUGsz8GtgvF4OCIYdZWQwdaiOtEWQiD/l/Rbuxh6yUo2lONTturzTNDaL
F0bf+utvWLdqlrdTYRsMbSBSGCnt9zW7nbmVSskXelWXmxT7z2Yv2h75qB59n604
uGrJK6O8m09zgM600GEgaftvReUHRe5pPDxiu7TApv/hCpsxKdokuSBWZaNBk2lX
OWvdt9kjLr6jAmzu/FGst+/PSOpZ0A51BZ4ijx97eE7MKus3nhEVV6Tai7bL6r38
L4CgMbF3G67syaA4C15V9/23g5MqhG+ay2e5zO9TajP4OowgQBkQ1XMwtBP6j7DA
sBFJX8tBSirGG3EtBnuffCiyJ0jXamECN9NgqxVQ17UrRHJQYwCIE8A3C6gOG8rN
G5XRqiuH4J+ESmM/eEHY4eNbH33N4XOYSvfrC7MlJ3KQ98sIb7ka7od+mQZ0QsQR
TgkiHindlG4o6d53n8xvLrLALTAiwzmlUSUZWEOyTx3wPbjkAN5No1NfUXUl5Kip
1M4r2MQ0H+UwuT71QX+68aKx3pOyIGPP/nc54CxTKkrGETDCT1vrq/C+P/UxHTbZ
oM1bK9/RIWr+ko1Ivo8kyhe4Xn50Q9KFz/xRNcSa4uTjx6KUlk8wY3DbNIAW64J2
kED43Uhvwcm4vHgrDTGL09tgZB3eKZTApENHxslqdZiMwejXHVL1/IhfF271Aoby
QY2+PpRpP1N6utIXJYX9hwQwQs6pq/nvgcd/1zI5n2NwhRuxedQvfC+ncFqKQ3hm
mgUg+YUvNnSAttxTRfArvd80LvGlrH4mo0lFG6yzOAfqoPsUXQ7bnOcScaHl0DkJ
3uBWenHBKmEsJSrBv5LTWAatfXoF1iPQSMGzzwHyHEFCAhTfkJ+cuFAtMPFyZcSC
DGHlK/nYEaL2MCaFDPMduks1lmvCFycbiUAlVQnFoNd70RzEWmdGUtSxqDh0V3j2
UfA3exLCKz9Nb4/QELaduO6jGVd5g7YiT9XflgF0N0f520es2E1tBTGNy+g1td8E
f3Y8ewTGJPTJ5L6Urvo7Y6odtb8vaAOYx7B/HnfTEQOZOMjD6UFTQbwM74TpTb6H
vwL7Upjp8YLsM31FjHJc9Rl1I3lxVyzTHhyx1wFtv9cipGVxclbdVjYrzLZIIZV7
6zaC3tZazkyFGe6mFS8wTZDZxwBGG/+8JVzoUGVovDpe1hnYSLuvRQr/EDyb2A8b
R7AQX6vBpFcRbrdRvDwQJvTXyuY3QzqJEC7d8qnMZwhm93lZJ9kMt22Vu6NZ4nsK
MuCiw+n1jkekyTMCLcBkAkACk4c58klt4cEour/dZ82j9Thntgd3NEJItXQvQpFm
i0RWWdyjTV6B1kLVQqsiB2a5J+aySZ+42TmKJp2Tb/tJuvTkOAAnNQ4g/+eBk8Zd
EgWleeoakK3/cToOaKEaQ6WnvxHHlFBugJ/CrZgNXfkJ/YgP0RX1bxzGSeloiztS
gUkUGGj9A7qUe7ZbbY9ZkLGKkxW1WjlIAmXGZn636JN3C4zyZq9b5sL19P2XI+uT
g+EtRFwy3qsOjj6R7nZ7pAZV++SNVyA7lc8f77ZinwLVbRC+oQz6dvsK4TVJLa/5
iXuDj2eEhY5HEfQPaMgKbxBEXN1pJ52eCw9Mu7ucN7G9arap+3EFeAvS+0bOZzTY
TaOdI896HujlLEprvafxtGH34M3dK1O7XCoLsuhiTNR8D5bjH0oregbo64s8SpFO
8j/mqUKqmdNswD2YLzSSAeCqANToO5my+JtCYlcNryATzPP+B12Qc9lF5lTxbDrx
FSN4uyFNEnX16TlwYI9f2rTDza1UE4BJbCbHzgXBB6iMlRx/WigrUdfrGwGrZudq
nIviO6J4X19uRFb/miSUTVfcibvOEZ3ncjUOXU586NLYVgVydn7oto5deNA6CMCk
AciYWa6KaG0YMQAJaAKEpkBVTLulqIG5bOPoJl0reits5T/W2i/MUNQ5aEuU6sI/
bSy8AUccNnvK+LbTMO61ee1njyyu9/czZb1uDAvQ/2/Ma46GRW6XPllpE5wBhJVI
oudTnm7tjJBIG9Y144+ICWnWIthzNG7PhoBksY43gaoVViBB+X0cr7b6luL+exAF
V1LlXnDQLzH1Uck/UNXvTtV5D3X25i4Bl4+Pt5apOspPa0A8XVvVIPXGgs0iitq6
yatbdOReyltDJ4iicYqAQJIj2eGgJ8GUx+8Kc9VJvNerE6Kqhev7a2Dn5PAPM7X+
BTOW/cSgnNWbDG+szci2jEdLfYudXE4LSurGCdnVUWkCoQ/hLB9KC2isBb5kwbhv
iao3Iga1jaP/TAuz4SL/An/OtbCPMBW1ZVdUiU97kZ6bi5/kJlbxuBPSESKF8o0C
ej5ZIXkym8ZvOdEPg3DCbcocMxp/IQQXGkum7H8W33J9FoahRVJoybR4WsjJn6g0
yiYZijAWSkwzJx2mK5GaCKxzBGW1CbrNvhAnpPth5m7titl/WLhPA+sI0V+Jl8Wz
Ko2iT6JZQcXgFprM2W4oBQMs64PtQ2XUPjDiix7sLEY12z05YYU69sr9H9jQcv+1
fx+2gm4B7QdGSHzQXxp5lZxm0bOoDAjarbfuw92gM9xrcXk9P0KyGXvgeAsUK44f
NLS39ZvsMtHjzhgbg7MfRxmu1G9NM/s3/Z/9PgNwFKrYbl+6nKsLIpS/ZaE+GzFs
Pe1fJEihJoP7E3U0CY2YP7ouGnSKw5i3JWFljbjstrMVsdP85x6O5Th8Pc6TcVzO
lJqq/mi4BiVQk9H1BsIH0GVo/pJVk2M84V1o2eH4Mr/sx21viP+GbQkl/z/wBuhc
WIur/H90g1D8rVapHFxwWkuu3VsmUMzVIeWCXCgi7XydoThwqOTTJJtbBOD/F5X8
S4SIJz+4kuK7LaSzlAhxTRqr3Pl18o2WxQzIFkSdd/IX4VVTB6dGS2ri6GigIRlA
se5rKBoNKILVEBME1E7ddEhV3wtIrh1coX5PB3dfimhZ63yl68JgRkFQQ6upaPTK
E1byJzgqBYSfsrjSNcKibcDaXG/LLzmYNt44rTJjopxuoLXic9V4hU/tUoSvBraf
sCI+ath5Rid7WDDd0eLJlgNRTpMorD+KGRBaPb9bV+uYbhqFFgC6kVSslZ8wuMFK
bm7dnQ1XufWxutzxtent/Es7u/EWGVRBaivEAS8guCslQGwv3myaBp4CpG9DaXyy
4AweyFJ43nix9qkd1PgZHEynY62cndPN7gh0Jgr/bthkE04mWv7WJr0dVZjWroTD
YoD6lJjmWgyiQhE1yf3DOSdn/TBBROA5QxZKx6p0PM5IXXj6BW3BKBjGf3LCBvkO
w129NB8ttFqXgblAebHQY3wRi+AWt7ne+pqj3TvVP+S1QlE4gXL1w6MKtRaORtcI
hU4QQVkqF5Zm0GDtl4Vv9sI3GzfxF5k81GaVqqsC4Qd1MiLUWkINzUSjkvVwIbyn
X1xhkPR9vWzU/Mo81TPcftwkrcNsSmLauiNLSovFCsawY5XekvCQchMT26LKnYYu
+go72Ll+h8BWXXEKlfYQE8DNuVYlHIPbTgv+kLjmERfVL+/HK55pZBcmtmQG+PiI
hQL7tyxhh7bDoDUzvNSHHnzmhCFV3drAyZ7TvGcDc5Z37eDRtVPGx/5ZW7QtBjfF
fKc6YrnTXrtl9B9wed3gxEHmQ9BB7UAeT1gwdZ9darM/iDaiRsVZ7yIhRABtXig6
Z4IOKF/C4JZJIPacaem6QQFpwvG9BfplAetxXfTClvsxkA8+r9SJthp46Q8f6HVx
E4/KnesAxz/ELWrH7xznXYHBpjhoc3W07iDXrAXJZidK5wdGpEzoNZZY6oGSFL0y
CFysBakLlqX2wanrzswasi0dP10KmDvqRJ4PdRRBadQke5XNZB+lOrq5jmb2JgOX
smf8yTyemsCM9exC74CnfXxTkjFraVsUGDnfduws8rZCkpPJaJG4T/O7uyXApv1c
1XwMyGkf89HWQPJ1lCCotf5qsoJfZ5CL+JDxwmg4eQRD2pGiEVcXGTS5ccfUg+07
0JLexY1LrB72QLSTfTR5RLMVl3DwJP79XTNTP0zjUfcwMcQ6IK4MhP/vWEXstgVH
PjXvG6tfLw1adzNYA5wFnBBNQqVZDGlWtco/q6qouP5jleeG34izr1MlLQq3kE03
/eOLFvsNrBeWb+56Xm49Hma1dwYvLJ9WoxXaJ4d6ZyvFuip4fW6p9F0MoeOZtEX6
a7mx3vQFx+CN0WJFGctsfZVs4q3FJJqA62WWUoopBPPtLIl3LzuypLYVpEejOoi9
BdkGJMviM3askVyejOZCdglShlLjPJ6xydOVQwB3rTik2XQAkRDNSnQ+A7HLvKXc
0nVMw24/rDnf8cgAkl83FJnQpzrTxuQoIoQilHfXRdUAgd4f8V146N1/pkhItxO5
zDE8KpO23hVnPuCHpmW3RTaansuv9EdXDi35TsX+BMdBqFoNEC3PeyrKEvt+KfWS
PYc4xvzricbJDo7DEaAwRg1k43eIMN+LVOCw8CIMspOfVZII+XuLwWh97D6Va+g0
/bvBRQ+/1eLherErGbqU+zyZ7k3h7Y2ZLbDINOvn27udmNTbFkIDQxB4y32PR1u5
SIeu+Iruo43giR1UXRdpERQWGjFGKTrRp9bt2sPyAgLStXk6AsJeH8/lm9M4d7+F
dHuNo1qJ2EflWQRHo0SxDCc7KgFtfjFdiKgEC4oLvVzrJAcA1qrsiCsTskDUmoBV
bZoTtm+An0qoCg6l2H/N7hdsf/Ym70glpzcm8Xbg5i6UuCELd1jSLZgXNqEynFYw
LqUc7R8OoTXBm8YpZQ83F9nFjV8mX3/f2786DZqMFlpeQ352wFyL93kkBNlyoHE9
gBb3oPgKLD5/+xqw0ERR2VQBJyMfRbhX01svYX1Y0S6eDqzcvglhd/S1MVlFmeq1
fZ9Q+s5f3muk2Fm9RfC1LzF8mg/J1xvbo5DFXZ7ThKLZiXvlNUgXCH6JL5uW0t8b
p7WpAmgsdjBZ4LzBgrX7/wMn/ipele5FYzYLwiXSkqkL6KqlJcwnfdmUldM3msIZ
dcrSCpks88GFZzSP9UyiluKUsCSiDON7dYXW/382BVuJcFCeJ1SRT4AeG+QNeFRg
FiA8tp9DaplvzlTR6R/LUvojDtE2Vf+fFU6yycAxLVzHOJha2OQRsZL4G4VqX2pr
lrm5e2SQGvyK9PViwtqclA2C2DbJBzLI62ToZ/LLOjlT1n0jrmpBRkY9+umCgrsy
7n/2p/aouFgY+vK1hsvRYpNqK8yqvXhmJNkOtL2s4w2+nwRWwplYwT/icpnPTxtf
mgHEy97X5ZCj0wAeV8ZAOAK682+2qGfxGOYA7k27tZwmCOCF78QvIrUSl8KEE2CC
UC1isvxtLrMdIoUiMmcYjkG6M11edsC39umZ3Opg0XycF6aOm+4uOCl1FHZ6PCc4
ZYSlppSYfqKPSwefyyeKBRPsuuEyD4miI1n3WAotYlQA6tjqn0zYTIkFP1AbBzr0
EpozsZU9lHIZE6i49No03oYNfk3fPR0E5w81lXsFraID2Zv+UqIZEcdcpqM032Ac
cOEjzleyepg6CD5/WKn3+AXLzUkqUhxlKt0zVBiCLNf+Moa+Wj5hqUDpn1k7A+Kv
8hu9B3hm0Bog1QIsNhbhRFbWyE+k84p5AQtvgtsXbB6TJP84NdvuEQxOJKTewEa+
krTlMMaiclFa+05C0l6zy2moojnXp027+7CVGsFqrV6i6VTpZh6Y7IQ+SukZ5bkc
CsynX6L0VsQvJxvFkC+HDDTV2vEeZN4XzobsnYII73sfDXFHzZZ5ucEULlkW8yDb
Dv8GLJxnR/lVbutZPaDB7UgLnXJuD+1J/OoLvoBT+eIYcrfpBWpY+jWfgrL0XOB7
OUpmUqfu7owoQRWfm8EmtznokrpYJN8Z7vpjvfNLvrzaFJFNncevkE/Xy80ZuoAG
M4cBH+2GJFNeW3E7FV1AAUfkk71Iz+b+JTnAyL20nUmuiKdkXTCOroM7Na3I5YoG
QW2ytmzoR/ipWaG8bryuKF6NhKKMbVOUqtUX3dJ0W1pHh3pUbeLoDxZdL/6MaRrS
AAy7TbysRob2+R8lS9IUygvSLcVSgspcE6R7tRHqnDWJv+L/YxO3Sm2HO5zf/WeJ
0SyvBChO9E9MqQxMwFkQxx5nsV8SYSVfwo87U9zMXNUOvNZMvcpc7zpxi4YOqrVa
BmJ8bDsrAbPSFPExmKXRANddXwyE8RVdQ2lMQcnukzNfg9y6iU7gsM+73sVs/Xn+
/+h7hS/IkkgG0jbOWnoeDiBrGug1f6B+OKEYe0ltp+0r6Pr6S5Ttez1jOgVlEkSC
uRTAHGL3ASfA8cpsYLFZw3BsrQEuk1S325TS7kkpo87zjnu6bm+VGPs4DyuuerSz
1dYdjBVED3b7DP9J11LHAN5tYgVNbW8avfH5mdax0aagrJOg7h+ZJOkgnVKEkW5W
EoE8G16CrGT/emkG+vnhcuepaqxH3OJ0DCeT5bFvlnpibmy5KGArWfKWUzgcnKJO
koqhcg5FlhusR5hE+7IlVdVW28VuUk+H1m8aQim5xRNmja08J1zQXaY2IV1apJbs
/PDI2ays2qYgHfRCOj9bVob9a/KwVjk7XEelORbhwNNOHRXMTr8rrDpCpbj/xCs2
1u2qDWE55SSbwtijiRGOBNX3VKKlmkimHW3oXwkgXPCax91DPSUMUeNBkyF2UGtc
NAragISyK0pAjEN1Wmr+1Lia0Al+vowe/pw7Eppxjc2Of4+WMtSk4A9NEgFfJ3Z7
y1zEykz81J/o3itjdotZCcydeKrLN4VLGA4KZOdzK0MmcIlIYu7U/FFLIrxyx5se
hDchlEn1NuORY8N2fWUTvJngng5pDjzJ2/p0jQvo1AG4PJ+xEvyESmDsZS38PSGw
V9+XDDG+pqN1iqYCfPKXq53tzc7/Zqoe+kNUFhSmT2moFlh6Qjvaf5Y+DOJ4QTWj
TKQbMT4mmmLsW408mozFWNabD9hkdIe6/AJL/IObi+XI8JUVL/F+YVRayA4NMwt5
aLKXjmZ2n1l+r4XOKft28Guo2LEAwU28AazTkQb4shIEA5y4b08yNYrzj1M8cHba
Z3DGqfqrb1mSVqU8d2nn45uB+uIJzIg65SqwTKYyR2YxcyoR5Xe9MdhnDSeiPa3+
N3FO/dYmYNQzXOSVON9Bh44WoPgMfC02XJFXgU1QSZLuvVCLnnNxU2tQAv9wCGcs
9bP/G+q7nY8nvTBa9OB4+CQ1+SXwpJJJ9EB0/D1GkFf2dtHEO875PhoOk1xNCa79
pBaEhYy/xtw4GIPNLuM0YxvoOjrLMVfJr9m+I0JRC/ovBeSvDtkeDK30/i2FuwOf
2H4uawZzaqbiQCS4lHGJsaJ37Ke+/xqHarqmV+7zl1aUP4wl8faSi1GX3B7vPj69
VX57CFearwekufGzBbbr5m0+hA9VZKPJx0s6WcBCIdNoILY4Gb91VMo06An06ATk
c7Fzm9/ohanBnoq8qFl1GgZ5tWSO59Av2/xg8yc8DsVLHoTYm/WjpE7YkyIDLX8b
7s7a16Fb7eN7emZ94TWDSXjELUIZd9adN38uiOfkq0tVQwlrXew8EwSwpkSdgcUD
D05M//zR6wdQ1T60aDoSpi7YwrXbWJoOkQ4Wnkfz0avLw0SXIgYTtECz8TgNT5ik
DsQrRQvc/j3tZHZIMBI9a2ISM8vyIzDp0WVSZtI6Vxs9PgabcAPlaYylXiT9Gkx0
LBMHvn/dQg/suhgls4SMUzy34TDyQ3n8iG2JrDpBBRwsSTYLZCEdFFNjr8/Wfk0C
1v+/Kn1tbFsOpCs7dDX7M5y7iNK97eax0hgcD/HtoVHxw7xWS5bbLOwUMDNu/SMD
tSuLi61aky/ZOyY9mwbAKR5Dzm0BfHK9RHnxWNJe9iWb/MAR4d6ogh6kBsA/tapb
oYM+QZh5bHQV1dbTlJ5kOlNK/0mhxpXb1tVfMrxcjpl1YZHY9SBvezylXZVSo9KB
x00RO6PCWCBMJe6xvOufcBqL2cvxJDtS1oxfHXp9RuS1WOIMqeacsw4ExU3D5VgG
8MDBeUIfWj5Exi0z+5/Z2bnksek+mayJW5LJtqv8kLE2FJVNoK4sn+1edCDUL3H9
+SgeOWF18sFmoFVQJbG4FZZIQFRGXXKI4pQHozfx4yKejFZ4Ehb0rzTT3yYtNrHF
zBSTXrKfU38QjeiU4ik8Nx47F2iqgUD2tMg4YaNI7Do8mM5gZSekVrG12vEhXPZL
dZiTbR+w0ad+dp/Tmk5fFhTG1lggrbTYoaYY+MHrBL5RCnBTi45nOYGNnGAJWX71
AfqKTXFeEAVAtAvW/SDF+ZAA2CNixRMVi09n1PCDA8PtCzFYRYMZ/F+mZBJBhB3F
ifYR3Uy0S8imsSHwPpT96Hig8duECxsf+zJ9jEq8/yndm95c6tc07uWaig285MsS
FyjIfzLoV+C/aRDPh++nqQf6JLXq94mx+QAMdm+1TJoIeMpcZQu1mOPx+1oQlhGd
vOe5MPFm1og+zYqnvA/6ObCaslwnjBnBntz/0nrCpNH/JDlMV5OOfMTNAcWXd2fG
w9m0rP3caEnAU8TJz8C6YbiyrVjU3QaOsdYCwzLtnQpIY+Oz4JIoO5DuNxKcIyJE
aQL7Jiqn5+DZIM6ksxiZuqJoMIpA+rMlVEcLggyzfztFsiBC3leYzGYqOk9byomJ
GowHFafvz4S9F2lzF0RyzvVV0PKNGm6N+Z+IIPXb7x30vfG63tZFlDCpPZ3bs3Br
YXrEIK9PBbefCSm9JGvYV1eJr0zTJ73U2VTtx99IYfNrp5IrImLSLblGNFfFw44v
FsWr0Xbj/5YXzEkqNQqjewM9QIMN2/EcE0e85UentYwS3sqW1TkfACglEo8HEfx5
7T9Ux5X/koIFN/SovpIQiS8T7wsSYLnlfKgf5IglapbTC5udTqTIxA1WP52Rg4J1
Jg+FWpr34JnFAB/Yltw9NvsTmXagAjG8WYPsZA4uwsRFxbo0/k90x5SA1yWE/C/M
yy/QGJWL/k7Wg8crlkj5cuK7hfc8NOONaAwSpHp7mgfpDn8UcsBf/PNGgcgfe8+B
CkFSJcyBQB3QPAa8SQUUiKoHSVyR23/ZCk2+EvJN8g2gKeAu3Idp161ftZTWUxot
vr8gOBFcuIAqi3UKW1MXYJ6Q5ZNwmHu2ZfNSnWtfYZQMqSz5umJl5FKQXsBCJend
Gc4HUYYGkqSujtKAdqVuU2OoffyF9d4NzLy/fmsGCx0doffbYiRqmzuwgr1YsRnV
9EYN7vjI3G8ZUTzLQhB1uLJ2M7u33E584b2OSrC5ziXZMOZ5q0SbeusW7mnI34Tb
8/JGF9470FmBtHi4wvjjrt4TsafT6Wu1fA2+7TqP9hYUVt0ShjsWoRonMbQGaKtD
NfdrBd/3thXLr+wmFZoV0b98DxL3D/U7ochFaZY7JbumIXgBUbCMTjhfawKGV1Oe
Aexfgk0e3lHASANdkvnj8YAygsWoauA6k/viM7Ub7cO+oJD1f4zV0w8rxoNRH805
neHKY1txWrCjk1FDKrkWVC8/SmVWTVD1WduvIsY6eha93IAi8wUDUlmdCaqBy7sL
qnUxy69AwwEXuTBa+/UvKW0g68kHQrQ/TG13efyYUMMQTCtVoh0K97DNWwm5UI0J
SHoczSXkoWKeQlwJ67GRNJX1X4ENZ0EPnTxZHdmzqrEus47KvowZRNmZMiWVmgpE
Z8Dpt0ZDwDWVftjtc6Y8oUoQP9sVhW1lBc534+4fcwGZdCFSAunWgH6GBaEbXJHj
cSXTIbtm1HhU7VqaOu90rr5Z2gT8ozhk8LR2u8ad1ZBcFn1BtKKjHZgnp056My4v
EWfqSr8TAKLi4J6ppfGFzqptSlSBQT1y/bmuJ71rdiaDK48m/8+xe+xbFxmVW0ES
432gs7cyTHMRjAmV3oz2NXMN27BYQ0zW/0fwRnYESKsMWq94K3sjxVYJwIaETQP5
yJWNLr78T4QuE43ph1Gbg1Q+uBwHlg40f95rECce0IfggYDaecS8rDw57Q9e19+J
tskCL2S85IRjYf+QkZm41Z/mutbUaSlw0z7uVtUhOkddpjJ/y5gsIYrzgflqDIT1
xdOTVDNj/QMJ+Dh2Xi3Cd/pS3k5y5jw0dK1+/yozFJE0XTlMzHL8omGZb3YYd1ik
DZKE68nZYzrx7tg7/b2foh8nWGaR5EqIP6LUbQA7H7/C1uS6nHm0b7cRjjJNUZEl
FM0fECfDkLVLBibOB1kxYvM4XGOe5Zah7KmS5B2RRNq1xnyC+oL87dW1WYCrGIn+
x/yAe21yhNCPBSDrykCgAQ1Upb0JA6oANPKvk6/Jo07Wn3d8ALcf9rgXOH95kAuW
qgvHwkSqp23LIwtjiyoLwVrFEmL0G2+W814fHz/+R585YzQccX3/2OxjIfzTFli1
Q6sSc6Hz+pDeZvn19fwuCAc6/ZCGQYYXSRsEvlOIyB6TsKf+KzSRznbMnzhiCldr
Q7FofxOGJNF/mE+yljljtVMUTiltrXH3PHqpcX5omivSbNY3TW98IuEnaM6vfhPL
dol8xLe/alqzbYui3mHIs6p+Q8TeQSY5bw4OGcJj4cQCL7IcW7AInwW2umuGyQcu
d3I76R+qMtO+04KUM5yGibPxk+E+EBZRXhSr7BuF8n6RVAQdnMIylA7xAB2T3rqJ
JaExphVaQ6i0qWrGVobPiyWRbgIBsnOFE9eB9klifVkSbCwU8xvRzr0MKutFn47O
A4teqJ/y++mFsYh04DcWC7b1udNNc/SW2xSG8En9om3xUtmdIVTXUVLFBamQfb0M
Lk+8C/Yhgf8XaKplr/vajqX1bzOSMYZRIE2T52iGKlOmNm3Ltp2BHjq7saIcpte9
7azE2kuFJ/enwfKTrvHqUhrbcZdo9ejhpVXswa41DL58dD4tUDyM7zXgZ/z922nF
KqqnYs0RfKBGGYwWqXULWSm8grKSM9PupS7QQ3oCipSqCbyz/C54IP/5m8u/JqG+
opZSjmIv2m6KSfnq0kmgBUxC8IJTBQkTiVCsov7y/qnrd9MT3iO0EBK/Bxb0SRvH
qk7Og6GR6yD6w+iERmoTUWnN4I2AZtIO1mEQtvQFC/1r+TCP2tJ9T4TfUdC9Bc3W
ttxmmjwaYk12YrxcZoq1pyGvbIIneOJCRjX52SYQya29bSm0hlT+1WfvGMK9+1Jg
9qyYjF16JuAdA6LfKYHZkkvPBX6pDwyDzDGmg4suvN0o7jd+xi+vhxEXVkaPJ5pL
G2hewOD2tiDR0xy6AQer9Xu96SMq5iq7qU4KfjBuJDC+7IXqzh0RfDIWQmwV3NlA
0rDuFhEg4syLhfTyU538oKe/BL1TItl+DvOcspDS+xHod9af4qxPJdQX+XoDzfy/
U2QXuvEoaoTBLW9Hs9T4+K7YjRJghA6sf8lcXQpZ87r0U6h8VIeQtxB06UPzidFS
u2GoFMw92iW8DY6yZLiO45C9kpkSloW1cr1bPStfsEfSzqgdnS7dJAP1fuciWY2M
Qc0AdCkLf1cmtjy+QG96gN7VpKgGmTf9GBPHIPKxPiCDtjcYuTq7JruNJX794gR6
nTBPGaVneBiouFDfMy6Fag72mxN6Txigngc/jIxndhNTjO5gxrSoDH6sJnYp4ECE
E1b6YDLUR47rRZl/fz36bqfmv+KxzlSAr+aRW6J2QLCGUNBy3hJjsyaSizfNuG/U
VlWkSqyc7xFzRlWiYkriazq3RRIJpHPOsGSRUCZ5Ob6B4my+4i40TCErPJN7HoON
2JNkk/ei8jTxxffxK1cj1oBesVlpKKb5DQHOPJLXQxRlSvFG010ljWNzYHZ/Mqb5
pyln2+iA6O0MO9WN1r6UfJuwfI+Qg6hn3Tc8tRRpcEiqKLVZ/x5ZbAXV2A9ms9o/
4na/Y5+NHlV5I6DI5t0vKAWSRwNbLaTNZzGwaSAjvIsuQXQbtL7wlV4uwCpyRh1l
QbXonY7Mk2xOGbYWtr+3jxEoKTmwANEfXVap3z+e09ZUyGNtQZq4z1N/8r9NWv3g
SdCvGvbC8sy3d86GY3hcfwGPJDW5jtxoJqzsZ7Xy5NOzw6BixkeSbEcaV4GWXCaE
nPAKkfhODMnqJW4qrtemYIxz1QLevT4YIajfTEP8oNe0qguPi+WSBo8yRcayJgG7
UZAlZ3VVwRapbai6OqeHTFop67MvYwq4Us+AE92fr8pn6DQW1QG9TJ4Hy3VfboyK
T5Oi6pJVJdEuGCmHjTLavdmyCRFDtpufmdxriJz4oAj+101uT4dO4x7UODf46SnG
RtNHZboxwy8RTMSi2OGtNAt5WDJdVrZOeeO1f2qdUXPu8N/heuxaO1Tx31ZOndHB
PzxqYjFQhfo2ec49vYdy+u2fEIy2Sd9r2fcJfz4YKUYAuC3igKVNfI8tacZnlhoF
bA/U0QRx+GCCT7d28EJ6yIEBD1TDEbhHIyMBstUVU6lwQr54ZWo0QtA9BUux4Xyw
8oVlA2XNOD0B1hkRfn4+zkjcVev5Z5eEDDmFBo8AYP0L13Q5At3UoIVucG5zN3e7
x9y/COgTQIY8ms1Rjr8YYyQZYgI7gcivVp3bQGzIbIpyry49UviT+9Pfaf9gRhPV
D4rleltaOJ/er7ycVPia5Z9/gg32yjcgn2j5D+GnL7f8XgdpvFoz59QwP/M95c8v
09+jSAiL/3/u3FaT4KuGC9OLaNieOVxlzqbX2TIVL3o/mjdOXWJKePRBLcvtt0Bl
pw8hqRx/dNz2FKxRT6Pad90SepQdQinUIgkPdymCuVccVbuttBa8pZ7laoJ5y362
w1BVsEPvZtvsXriWCLYvIgLqXkSJSXvEC8PrV5RnM86KttZeWqdyK/mTH6A59JhI
aEEJcGVsns3tf1bQiWvg2ggsy22s0nAK4Agx+uyR8dqBvqGPd91By9+7NWMyD8wn
XddME8u6SZ5KwCxvrkuQdp49U36kwvNjHrMi9zwV13oQ7LBt2Og8UiZOHwH2nb8L
Joayvmq0R/W29ZTgtfE8iQqusA6O3bfsejs24vNpMZLMKtwvE7UxYiXU2cVxeC1H
yN4v6eBfzE1EaZXcPdlJ04ME37L2TGQzcE6KPb1dZBltxFeNQH1em7bjXnschFxy
85YpA9PwPhrR/J0+tSGta3FcXHUypato8HSAU0//BHGMlU9JtsMfPq3hJM+8ACxR
6GxwDZni+QFtURN3C1axVYhSdYBOkHtMNCxnf+7qO+p8FleuG2JbbZSkeKCc+nSL
hBjcQupQiSFPxbPKrdxerYO6WcT6sRkNUyvVpThxH72ZXbJKAen9OrTPlXvoLD7T
4iin9+Jn605WQp3G2TB1oVig9eWnWsOZRPdbiiPnmeoJJ92FdeX3393oTruqS+8f
jNBoY+QEJR09u+BkGgmoPO//YfmqUZ02zFFGJxlj8PB2iTUaHz4ybMOH61e3sX2z
Ob6lznC8fkslLJm0IzZJVzERrbB3Er3UHn2QfCR0Ql3VUgPhtdrYFUoD7ufQDFAR
8AUHphAqLhwM9+6VBBz7DVDf41UPBk2/Q5Si1HSig7vEHryLgF1GijSfbs6Z/9hV
xTX5l88tuxQEJZaV1ID+y+eP5cOpZigngW4OseQkpV4mddaDLZGS6aANNIB9Nuow
HKMWiaUTwphtZHI8nhnS5upSVpRaN7ajL1YFo2RzWu44S0jngR0v1ZQcttWjr000
FkcMasrbsAINT/eTCJCj9CGR12OerHoFnycLwQPVSguEvGJNei5ZVk9hkz6Fkeuz
vCyLRNCBsXs2ha361FdIecBCc3QpcauvSyQtH1kwIUOVkH0Rs3Y4U0wUPkPEUG5U
EJQmhOyhmBqXb4bk67UR9eQ/dspfEAZuhP5W032Wg/iXGNP74xZrHydmdmWVWj1F
gncsbmHh1TERbnqg1wfqEhGJucjUHM+PPKqhpSkThZr5TxudofUZscqR0u/tBxyi
MjfRZzyZARNboKtQHDFW8XbpmG3Ky82HVNP98fU65LbpHsBbLYbGhoaL9TGaJvam
mYOhdzaQWESwAknkI+VKfJ3FPVVa8h2yOJnucBum0+pbS9JybBQhgLIQVlNtCn6K
RdrfqQJDxB1bJKdR6QX9+nIVuZ2zhMpws1zX4sGByxjk2G8/ecom+Ho60MAlQHqp
IFDy6IFuq4j0Q5krWX/u1ZlfAX+pMcLiITFtlVYKaHJmu772Y2Ar30sEpVYvdZqa
QVTvFQeHXPrlUwK2OnZPENx0FNpkRDlvrE45Mu719z5xGpcRTP5QC/JQ5ZPQEmyl
53PWS8BVKPdUN4kwwLHv9Ic70FeRTCy4WnvZjwswjed3F9q5IHNoVBBlXN6zlXP/
IXMrnigk9k6SIRn1FIWualEJDhwjmct9WuDOvwIHAX8JibkHwcJ11slN1HfuZBig
cK0CFjL9yFUb/2qreBdpZZonm7MDIN0cwfRDgH15D4JbFev+ifcBcGilxIRiD5Fp
GhZZHlaDKha23SE3WAfk8CScfEJMoStlGwRwMfipFkYMDFwOUgi/JpRH+fzWR+FM
pdVsYZd/V41PMp/8y4nPijPMjOhK4FM0ZdaiJ2lQVwhWAURw8+rV1MFHT3pllOXh
3Qg0liApR/GD7D+fKQeapFeu5TXVgp9ixQdLIFHUjIz05AyfT4euHcZW2IfXeAKZ
JgVSU9LZO8t9+0OnDIfZgALm9A5P7gPEgWjcwrSYGhOPmElWvzRB2KTRiH2AtXtJ
xg1l6acHn8ZrDPcqKNydQCkCeS265BiTSOT2k+L/P8BP8uyiLGliRDoQ0yzIgrAO
kf8BeHZ/cgGa4nG6YvUB2iMHFo0zB8N2I4fa4pLTHf49slPST0pOFdssTd2OFUOp
X1v9ktmuZ0mf0lexhbeE4ripacmjIOT00hNjslwDg5KI2lCO/sZzIkDhQCziHlgT
/gVYw/fhRL3lUxU+22rTY7qK4yqSCD7kYMdwa1z5wM8mvU1EBiXOcuZlhtSVtB9v
fLFjDBHlkBieGFrrDWtYbgp7Wr7vLLulKO2VHAx/qJB/QWqI3LAhBFRbp6dBmS5f
9bDUAGJofWtd1tLhbcSXRR+zzo8IVeMfi7DevvXGbJBMVfdgjabpXIl08s/m3kru
31OmF5p1zEVroePPFyo59zfSH9GJghtEAps+omu8zQQUqd/fJ09gG0LAbUPlcmYM
5I/t5Ho+0AKLYXLatKyKDmNMQIdRDCIGSlL7IbxrlvJXst/gRdvQKY/pnr23OZTl
hqDTE6JN96O+Nw/w1H61VEwNVYOJKC4WTP5oVHfrdQnPG6BuYH2PDmm5fQoIZyJW
EDvqD2+mNee06NL2qvOtW/V/mZ+RQJwl6FVRbwK6ijxS4gNrFPBtcoDwcqI4Qfo1
wmzEsYOXnT2DQFItngindQ3J+ZQsStEyZObHgzuYGTLVbyc1lS/xCYZsmmHD8BD+
CutkHW98YkVXQTOsK/xRVwg0IBxTbGriPD1qFROmMgRmCXAFaBBUS3FOxI4e8Qzq
qxtnjiUIW/Bc3byU1aEJBi+FjcyrLrUu7FtyN9L+RnvFGx7wKoZHpXW1gyXbmcUF
xYgdFlyr/Ali3W1+Qo6+3IWMuWB5DPhB+cgXgMVL/b7E3wNcXj8baqDs8GEEobTb
58nEdlaeyeaGc1joODHWhQd41hDjf7xbwuziD/o5C+FuHUmmgTOvRLj79o6pxJSu
xBAPDaCrQrI4df7g5pkqSdbRR3fLq9/lKJNJBpfojPBMI5dz1a2KZrxXKKOPBue6
HgUcb8CpxFOg7UJ/1aU9rWI6v2SIg1Bvipw138zoO/EqLUdbW3Ews3aOiRyx0W/3
FDys0QzmWCyiA6Wv4ZH+XphCmmNshKfHygbcH/CeXcJz/XuDIq9D+k0Mk3IPvt+y
D+s6h4ttrUNm3rkx+c9SuV5dAreyW4TZPkzMR7Wa6RP9IVnOsKxsLWCcdjE7r5f7
9fnA+eksWpC+jA869sWMPAFopNHqAKBdyw4hcADv1kwG9Lxh6x9/5zFWoWXeb2ho
fpkqzNFliKES3zaOz6wyuD8/DGKpmPmtD5vInc8mkJvK9QZyD/f+ONnZiOjTQAnr
mRvvsQ8JpcXDYA0tr/wEQ5fdVXIqkoqv5dfJxkRKr8qSWbrBrpQ6kxGl52ZPJwFL
X9vmHQx3EMJKayRSeagEMmePb6JdFc98zHEJcXxzo902ZwKKHkrmJ5BsCTKNkTR7
w1tXvz/OcTcdqbRc474seHBArYKQWGQ2h8whmJQwNRrL+kskkjlpE6RMpiYTiTWu
h0BRAQxIA7VaY9gP1jkQqvcxHeIQ/O4d7rrKi+jzP+7jWVIqiy3FbmacXdsFBh6d
mvf5IdlxrUSCEPldJ8xQ9nEQ1AZULNsEQF/LvuGHP8SMXuQRXLxM+8VfNE1SjVd3
yWkHoOZynLbifxCHn9fnPKcUSJn9NTWgsTa6FMustUpabH95fywq/qRif3+7jg8V
/Y4ej1iIeg1H2Jn67OLK805j2/sJewLPwan5iPotQRuuICwY/Vi+BNIl4tpuWPIH
466opEUUazI77nuyBui6loFy/YuzV11inYgKQYChTNktNdYLEAQTCd7rc9XV4PmF
bAm6OB6O0PxffcMlkSW82yMVito8CO0j9ML9px8+5zltBgjJKwgsWdBzTlnB/6PT
MFonN6bh3ShH6DW97HxXS9E29JxpBb3eC1E07TKeIOPelUMzMuS029Nr+UFyKon0
DFQxJgsAZeoMi5os3FC3pWG4ZPSp8AtSB9mp5cqB1kaptSUlnN+krufp+N+G7hSd
wREss+3F0pFagmgatLcEEXdp59RLyPOeHt6Zl5yn/KIJG4lKbjdwb8+/vp8FkTAB
lqAjC92pjB96p+ChpmDfqK8LNm+ek8uEFLsTKnNNUYtZsg4O9cDrM5ZLwTpdZfsz
SqyJ1mi1J5XLa9fKq6uzvjZgpdaWa93Sir+ckhzwPGKSib4X2/DVCaF5rPX+FDDO
vECpsZ4GefoTOJBDzJW6VzaIRZEChPlCLee5HNRLuoLp4Hb8fXqrnCPtjMPxVda6
wL7h267vCslhYh+pT4mEXUkA+r8ARfcrL6MTAN2YPBvQDoF8z2bPyb1M2P32W0gV
r3M/Y6lxVubXoFMJN9eRpH/SwIKEDsqv1zBJiyVFod1iqK2WODCspyl+mPoJNYHx
jbaiTlROa0H3MjfbeHGjVxpX9/MkJDYGjc54tE40WgWXmTsPhNxZtqahqSWo0ENE
yrzAWcbf8Gyww+/TJ4BbD0RVZ0eUWbK8YJZaOw00MmcR+rCCSCgsRGR8sDAJ9C36
ycRpJQ8M6xl2IoySgnsmj3K+lmWjf56SyMmzzdqh/NfHX0jsrQ2XuBayWMDYGpoP
o+R7KI9J+7VXDG63/gznOWXNEK+zPcXo7yJ/cL/LEsjngrJJAYknxhqbWT4fqcbo
zG6qLT1YlEkaSWKVFHX8zpPgis0SmpkWbMxcg8+oj/O84UHUi80BcoqMWuGEiF0L
xw5rNmciQ5R3m12dsPIhIT+dz++YpfnmuxgrX5mVeeXwNxIXvaI8tmT3oHvpY/ls
LvMyQlVkNRSO/RsN0L3dgvsCZ7T2n0PNkEPELlD0ia7uQEJmuuTweleNlvZHzNCX
UmxmrYRbn12B4OwSt9wnwaw8Mg4F6peiLruR3VDpNmoo6Yc2dFlBcM9VUOTOK0hp
MFHR2GzbBrNHZDNK0Q/khPLkb4w8e4pn3qThlxqXcrDWcqip1R7zo9pSciZJ1Diq
MG62BTOlHNSOj5q1DbVhrTDUbP6oCHNsQyKPGE+MMKMCofmgWad0p7aaUTGVW1pX
KUEcxNWpobL+ARzWxuwDi1onbhg1bwomEAFe9xsZDU5hG6o4iWVLa7U54IVi3q5A
gExnLDh7mjdY3l4HJRHEGUUebK1Gt+aRl0xhcT/9Jsz0lxgI/ZX0MhNPKXhQTjad
UjualhcDMHt59uv5NVHs+ZCueBB8Q6scLQpGOKD9anDty3MWzoR6eqzWNTuUEjF8
rppB9ay5ueFm8d3A08HhItIWvJJhjM0R3ueZL1uIDfDHIe7CH/iR3iztPojrwwkC
uKpuaZPTzeAXDQR+XNjwh1kPNNmEjQQzPYDuEmv+/V7G8UcLebmuaMQ3NboG0M0C
bS0r5vNnb3Zl/pRHckAlbU3fJivLmrAx24nuWJ2wpsfdarHTz9OrhRYoCyuRWD5L
pmdo2iRGODk4km5Jo5dwZebu5vH0f85+fdzrx7og6dQaUMS/Cm7kKE6TPUBzceKy
F3xZyb6oBk0Se2DGG1DK5mjBicbYvJF4/yKXIrT+LG9y2i8GBMv82Z3nR2wMBJ3k
J6yUluHjJSMZCWKxfmjK5EuCAyNGlXTNl78quTp0/zOqKD4ZYunc/Yrc92FMFtcJ
n8m2Jzu+MFfIkzqkm2pxI71IVfGROfldAXImX2VNWvtZ5qEXp1OZ/tag9itT0wXG
n0CgR+6+TGcL6KHNZYehpzrmVdaCFJT8WlmPNOrAc1QgNuIRsGWvk2CfC339151n
fPeAXTn5TOCkaK0Lb3ErFbWI2itFUakjuvXmlB1Jn+wZDJsrG+8GeEIjNOchYTki
2grtUH9AEZqod32yhZtVFwdQOJTUjKkAZgJmVGZ68p6dkJKb5tGJOY/g7mH4bnVf
aj8uynYhqsrNoRn0xEL9X06Ok7hcRunN9Fj2zRHXuO0YCRZ5p3KN9w9KouRfEVOj
E+TOIu9RNnQC4Kn9UVR8pfVWA1CeIPD9rX3/f0DlVV6wkyK8BJ513eljM1N1AMlA
kKoW5gva5EJzbZgXTmj5BFh4J9giIDxY7eqEav2K516SfKLG0Xne6LCkSDiienTg
4ukcnT2efOLI1zyxyxMTkdPhM9EFe6MVGGZHPFLpvJyy+S/qUK/+wqTbLFTLImy6
yA2eqO1qVCb/GjQf2PqsrSmVvhaY7/8AG8T//kp0UiJB0u09z+2OPCUzNDaCpb8f
Tiix8FHzBgQobEN8vcroEODgH/VcBcK4U8bnzZwscRODrK5I+ea8InR7t/wkeqcO
SWQs6mDMY2LKGYEA/2ZB8bcla71UQ1Icf8cA/Bh0ptD571nSio9dGTaAH2zEedC3
UFiPuYIF144CNTd/gDc6IlX7y8E0neYwZrDwg9EXPZ1tTNwh9bLDbiC3iVK/rn3A
5/dmYwbHJxHlZVDQWXweqZ05BJ0maNHQ7MEHpyFsGpUGCdey7zP+0fUQ2XXqo4f+
TykhqK+QTWQp40Z+/JyDkZPxXoXNS+kj4dO2M9B2PcwcJQfT6oIc5dxUQLkFgq26
/u3KzigJMisLD3HFO+6uGY7AcuQPPZOBhYIuxXwzFjLuER5nkwj19yeCLvpztGAw
m5FoT68Pn0htHYmEHQ12Mk87/9BaoU/D1RreB1JTgqPY8qVvFO8PNz8kQ9M9PUaV
cAyoA5yu+zBD76KOFrPmpotiAYDoXXiURDW6F9Qv25Hg8yZVA4dvJGwBjATBvSml
scfWjAXrOsYNAWSrkKrRTgxpYmM3t40XY0ItYS72V3kzAwJVoiHZ0vcDj92TF/aN
P94dPyIRYBUXG6gr9WlzOxozzgrp9qhMou4F1Oe0rAhiIj6eo1edMx8WYp4YOvpz
TMBcxp0E6YLC0AXMLKrfWI+KGVpgCvMHMcQAiE+3WLTXOnAAlxnXq46JZ/6u28VQ
RYUEr4YoD/KlultF9UhzdNwDwYjtyYfgysu84VHoFeQYQ5oSM6Zf/TWUlstR2kVV
w0nTrmcHRUl2a1fe0UITu+YjFtQOd5lYiaafHb0S7ob7xEim44CCnC+O80LG17+v
ZT0SmYv+z/BuJNItv86mnmEUnrMBM4mZ6OBd4ipoL8fM3FwN3MmzpYj9bHhzDo8k
EPRpCtSYmFIMOt7M5OSKTUkqPtNv/dLcrmICR5l5lva4GaWvCkm5euaO7YmtnVZo
Q+9vRSzrQLpWou2SgyxJI+SXJlXEqohyN7dN4u9CppAlapPiKV+WFo+G9OQONTEP
LQhacLQ6H2gBSGq/o+GtFGsMIEjvrnu7W8ISNm5xKTPMhsz6GTBiE4xK0UqM22yo
r86ee58nl+cG0f2Xv76v1fNlWoOLS7bHNDDT1FYNTJTVMZ8t9jZuQ8LuCAjm3J8f
9zdSFhEg3MV5WUo786v2Xsmachl8ShCOdHWA05GTrqbm+OxVUYk8iurlH+4YU5Re
aFqT4hQxaDBwNE4pTn2xL3yGCPKpJvrv0fyWZFDkIaBCsGPqNarG/ByhnY85KiQa
CO+cHmCI67l1fL4spCrUUs+NJbs6j0ccxyUAlvvC2BRKdXMO5YflA46yOHjkGDqL
kFrhKxgw2Dl6La4CCmkED4KzzCjS/kEV2psI+YNLzQ22QAhXicGltkLrhJ0JLYqg
6ZmH0ul0hH8L0k1DyG3oP8AWmx0ckJ7yFUq9V8FIAmLY/cKvJy1q7THqsHLrQx5D
naCv2VhnJSeCFeKZH+5QCg3g3n2W/ueH1KoQm9BytWVtJDYh+CJQS/UzZkyuwyFr
ChzNwV8bxxIXyM1XA6ylOzhJHXgJmQ5lBeC1IUwjPlSgREUShCh6pkWkleL2f+zR
hLWF9ZhYynLdQN7tH7NtPNjISqEvIhlmBluKae4qslWL8x4qliLuS815QoDyAKTU
sQYwJsWHDn9kMkk4EuwBxw/YFY1NUm/FzjzzE/T6E8L0PWozJx/HWgwJ5SxUc8kZ
zggeU0JjW09Rb7s0HfJOA5iI5UnC72X31qBnCUmnpv6vmZFF3oMMWzmuKPBgrcDX
5ZpduETQZ9gw+aUeDg+T4RRwFXhIMPrKWJVFOzbhdH7hzvKU21zu5cCn+yN3semr
yVvXHsjqSxmNwxmZSjPTIhb7TIUHAKOIfA84mgqMNSDFA5YUTrGMU6Yu5v2ks3p0
iJy3DQOHZ5Ax+5evegUnszMLv5h3RhpQfy1Y0Tyd72XOYGi3oRwl84IDE9Ivx9Lz
a+kpt3dpQ3tO+ChaRT2dEj526iPZGf29QBJfMes+L877zibSiSIDtcEERqtg4Nr3
0QNkP/VeOLUDy/QeSgT81TT8fDeIozy0iiO+tgqg+/BXkAiLQaeTQBoTPUFUDdqF
nMGWesWVLLTTbRo3HQTGJdUJMS3yBZgW9UI1zbC+5uqWhDmIgFEp+8b8t861EtRe
oxYcZEHx9cZgsjZV60s+zYtsKiNO3E+djsPadephePYFozuw5oTNu90GH0ILS0Ip
iYqwQg0yYlkw4SAh7C76iE8BTkHG+E6Kg8Vw60ZCnNODM6exz1b0V1om/YWRmWzD
yZwF3IU2jAnBPwobWjAT74k+AkBhLcCtGxEp0K+lEUC7Y1+ctbrmE9eYlnNZf4SG
r9rIjG0ivedDcQYSGZkFldDXDY3HZug9fdAnoCSgaupY5TWBe+MQGzZl+xE26ljw
ikjqhvGdYjOA15Nwa1oSfGo9C3Du4C3lOx8B2E4+2nZA/DKM5gKVrLurwDnW4PU8
gHYkLFo60FvsCHc44YawyX4MV0WObSs8qR97AHI82eu70WUm+NW7NQWzuUo9LU7v
C7mhEW1EsRsQNudywh4gL2jtzfdpJzxxkqaYcUlpx1Kj/9OmXyZEIlT2/OrDUljR
9+rv69FknV96UUi1q6YIiBY3UrrmKdCAJuWo68HMhuUkLgCxE2U63SvmZwfryrYj
B+ugWfsdfrmWs9JVzc5j76HFFYVz6g87M+JP9/PnBB9vVb3Q/fzf5GkzSbgcKJr3
puNg5xaL3/hVCsZoEcjjTA9l8XWXM2kZmnyYR1r+hP4boCHeTZMSYI2vN+ORNh6T
HndetyoMEq5KGj3k2hsEhHfbn7nQcyYD11AiBH8/KhZnFGthkHto27SlMDBi0wQa
06bD66caRqYkBYB9qh9ZF8WaunKN6QHsqLomG+2rx3/6Yia+NUgHZPS3PsAW8tib
eWXkeZ0h3RhF7I9UHD5GWeE3cfywKxF1oqrK0Uf+lZpagg4hO/YbwYea6Dr2E+i9
gH6VZWolWqdWHNxMRCcGBfQzTxHnPwMdikQjxCro5kOXDv2DKbYKRVpuuImxLKMR
W6htKr2hVBE1/0b2vvexmMl7x/nN1N0NPkWEaJOqRpPviNoVK1cDj3btfnop4LUo
erne4VyDOpfsm9j3h0lAXtnx33tLJThDN6AIVnctxcBThyr4rS7FHI/P+ZvuGwSg
RrjRyvvcsfe7SZQTTR9Qv+Mkj9jOlJOAWbgBW9DYEfzs2OkY/5F/PBgxs5IAWbj6
Pvc5/kAya4CRsMZpWkk4vegqk6sHLpAOYP3Z86C/g75olSZn1WKsRn+qehgCD515
Hu8uAKQYPpwJPUAGoRrlY/R1tyxTRkLqZ0Qs/MTxQbuNvpuHBvag4GLoOuJ2IG5R
mgSV+enetxvuJBy90vmBPSdWbXYDQrBdwrncR2uMFQ90tSu3ao8mtwpJ9Js3gg+E
NOURTK664P3Yem0oID7QLMxLwxzHLSBWxdbGemddnPOoJN01QmE6VOFJiRCwz5GY
5DdzoIlQLUqt4CLaG/SbDsOFg/No3VZOdfi/q4zJvwALv/VPRGqvK8GLfHziuFeu
r1JaUVN2Uxr/ajPmZC9Ld0QP/4Sk1AloRH+C4v3dVjBh22BQpzNZ3aHh6WnANOAf
zwX9uzdH1Spgy7rN8PnLsBrMrVoFnS1OfaFhv4nw+LOoyvRoZOOqbCjpEeklUb8p
JZZi//Wx36VOCuIWSLCp2D9RWJK8IZ/2Fv39iJOR3WPE/VIRChggw+cznIbu8wF6
7jCDSwe+ztf3gIjde24Wn1aHpdAhqZORYWW/caTnPW0WXNB07zdgVX5wtFHOAuR2
UvbLId5FUN71IxB6/Y6ZgNC8sVMTyvDLfadoqZO2/SXvDT7cez8rbUKoDUHIyrCL
+qxXBjj5WPApiFXaCz/XI1P+0LOUxnEaPegEzYlLRyURDFotaukPkYZBifVWtENe
Wg5w/TdFBz5N2TOkMn+FAPhTk9eUGpISxjAZe53z29f6s5MHexYUdlFaB2ZtwQXU
PfJ+HVeRAk1URM1ZYEoCFaOnQg80sk9A4JQB9rkdMyH6WW4hODCqgGPKJ5NSVCEa
3Zd1xP4cBND4pYyVmiVndSKwLki8gc/uzGJGovhHBECaF8LfeLNyxJpUxMbKFOKF
6hqtWRKSe5+JRdDCsDzw+X/WL/VF++Bajoz6FF60Bic09phhBDJ4PN0Vpuu8oxXi
y4LmaU4LnHuKYCPVKAlwEFj931kB3OB4aWmi5VGNGtrchCPoPZX3PHHNVjdhCV1n
Djc3xMEwgCPI7acT6CaB42a6iUboKVaD83yhyXOQqnMgSYt1hLG796bx4MC1w3hM
YSkbcpsNb1ZNC7eMunyNKm0Z1Nh/u8t9qTCfyn9CKMu56E7yFgffEZobuEkhAy6e
6HNSfpSEruZmHqobg9+0d/ZKu44/TrG5WER/8zvfFY7LfYsNC/QdBdy2lrAQ6L2d
7UxA+yFaYuIZouf92GIteHQ9WIT7ytUPSiDgF6vUNkFgsihzJkb6qntR5ikLIxSg
TSLy1VM1A+XTkzmmLv6EWU0flBqFTegIHTt5DMxlvo+qYzD6J/vqesFZFJ/qAzxC
Omi1UVhqITKuz+KOXLeYRepT5+GnS2QoPSCDF7GVEKQig0ltDbHxQpgrh7P1tbcs
SqxRofvt0an+a03/dxNY8iXzTktvJ0zSx+2qg7ikQCCGVklNFokjWmHRGIwx7Cdx
LrqOftqpwGxK7djMdmnn4wLAMJTNYQDNgnV1E7A+edp2jnd+JMkipXg7zX1PpwJf
Boq6IjTeEcEgFGi6mxCUv/gOmpXU4SigwLjAsuc1+s0gcqYSB8mHeuI26gOWs7bv
EO4sbdRueSB+OF0+ybZU6dzn22kE0bAYoswHYvWDIVwBm9ddW/Jau7ELA1eocKWM
QCZviytN9CeyoLj+7myNaLlnoj7nirhbllFMApYmV08TqOVr2a4d0zUYqAIkQEsA
kHWA3vZuUGwB28Ux3pHXnWvXoFSetzbFzNEK6D5Ugw4YyeXYbno1Dx98k1BA1rri
X3maizAIDDefbRiCzmKspgb7nIywr6jo64srUyfw6eatNDq8ow0Phw1vdO7boNAs
ml4F9I27SCJRU4WYpSCdW3A5E8OXsvZk28ywfQXykIEieAeZN2YoJD8BPW+Lntts
P7rA5ClSgS71si+YYdoeub0031IrkCCDyo3g0LjkonQK6fUqAp8lwDGW9WsOx+zU
tuN5Ci6X6J8OZYbjWioqp0/7VeEYQeBX5MHxAhBVXj6thvBCi6181Sfwg3xukq4R
oH257/UD7HArcWYE1A9wKmvXoV+/wv1ooLn2xdJsMqEV3sjD6atgU0Vc1PqoERZz
klcHGGbfdIzbjCzcY1QxVeuxe4oXdkiJXweZgSu7xQ57iXMIFqVurwgWtj2b3jRu
xV6gxInw6zzWk77hT0I1lheY79jspElx+Y5tZ7/zhClvf2RXhZXFqEtxd7LKgTkp
vR0Oc9paa3EoVYZLRk+cj/OCvAAbj3h/CEVpllNLjFa14bW8iqjs1ixeR3di/wEq
4kYNLIBoAek+9XSVoQ4DOlRqeD+/bk502V6QJqtvf2Q/ZbP8x/CwSmFjZPxQAGOl
XHHgCCFrGvf1jYiKlK2aBSRi2GU7JRw3wLz5YxLLrto0M+vHmMJQz3tT6YukASCi
EMLoJPwNxVI8xExwDHrRDpTeQtUFRF6oDpsYlA9bR3vCx14CZoffEeEPGkYFb8Vj
8UwJts0A077H/ATssy3EaFlm80MVfTZz6Su26a7Z6BuVNMjrtPULflZi617CtgAS
do+WDJpU+4WPL3Yg78EdC43AKklFGuMo6QaM5oowJithxku8DpuYE04aramvp2mX
ce5iueYXYRhRoVEjjSCuaOCioh9Fso6QbJWFv54jR64Jd6/UqTONDgGRjfoBNqsA
iKAp+qdMAItrW8keQmCvb6DgBZM2R1Wm4hbX5pxC73YKU76wmPXCE73adVi+jBJ/
NZnZVpLR0yg34IuGm2Xn/rdulnSKAc24OPCKvSObM7A5zuryJVELv5OWc1gTO6Uo
BgC0vYAbCTzGuPKiH+EZHZ6k9B4u8dpOnBYcACtSiafYsSpNnMmTVR34PcpDOZwJ
J4Ug4kuv5fFvSfGk0dBCRcNEUSoUDSWa6xOpAmmrVhh8KAxh1UfVLJNoI/XOTKVv
HwcG8HHG1Fc7uLvJQvM7imVfZ5Dy7Y15fkQUi+mXj9RMoJxYW6erEI5E6oU7DSem
K7I91McTsSjTt0iPbrjxd/gw2oBsJHFIGIpEOC/Pft9MYFn6h1XQWIrK7+FSsmW8
tOODJQH0QdWk0MUVkEY6lyBqdPWtlhcE9N9I15T9x7EB9txkrIKXB/CiFonwxL9K
lyR/eE76EeBG3akETabJLttrPYWSkL5UEhnGxAlZ4fX65B5E4Vuu5yPYrI7MToMG
OWjLo/pu1Jw4dbqzx+vEKtPy1o8nKy7MwHp5ssJ/ePwuQgY6s8zJPIWDukPJnvBa
p2vcg/yKEiJmqsvidn1wHh9qVr6+3MfQuAx47Ts9U7bVNIki41+AD0SiSyf2XQrr
voHDDBRjaQJ/CkT57Cc/gJtXZKQVSLpdGvPU6h1dUkXanp0dBuhPVK7E0xAyPzVP
eXB8bH8SCy2wihdEBq39Pt4G33HhgkkuuNs09h1QrOUzhjt04nEbZNUUbnYKkeXo
m1+Y4Wt0MEK5iB4oJh622SWG2LtxsDiiYVHToUnkHGQpx/7ifAKl45Nut9qCzFF/
4cgDiDYlbtZQ1KV/56O/FbOy2mgh9QGAsQgA21RNYTIy1YL136cqZzco/qxypTF3
2yD67ssMLpB/Mhe/E2F6oj4cyVt01ho0LrDVj6BuNCvX6WNBrSCZdkoKr+fTXxUR
LHV4VdHO8WtxI81XuxMADzdOdMRmCXxsYXsuqR2UUZlriZPIaFwLlIAoUeUTOQEx
VQrpNTv5RILiap0OyVT2g3BJO0F/TrtaPER5n+z7we5Yvgw0y5UllddSOzo4WWsA
e3A26s7mha9OCpLcK8Eskp9gSBi/NXIqrOfG4dc7VPNdw0wqIqUvxXa9YGVmSo17
I3PlcZi1tTq1uLiexFL5yq9HN9njC/5dXMsQ20PjJNTsanbImmeHsOBWN+mixW0X
BVOd4eAOQ3Tagu5CgeM3GMQHRt05adLgooitkybJBc+C0YZwEIE28te0IiD1Y+88
6P7zGklDx+6fK6VpJ96bRJUhh36LkSU6n7l8FarASMrwtj4h9txeVAFy4lz6YDH3
oiBoUEh4BTiRz+ZxgLCpB+NEbekVrq/FvFQoul6AlLjcgCXg0ANRAPSMbkgnD42/
yDSmxKR0mkk7RXIwaB8+RgjBsI8l+S+SYqBFGKzPxfYhM+3AkxvClrxXSvVrQozN
wBZ2Ivc8//bGiUuDE2syMHTwakl4e7h/k2rygHJYJrVRCORndW+sgvZoYgEZ1j1t
p6KzPxwCoGtyBheB1O84j4JS7Lm8qBBhxSa8ABJhjxP52Gnmx3lwJxp8YUG+5APU
SdzOv/b7NSA4yvTrJhpQepLa3+h7UTd5VViBZv+YiwvzAUdP755LSJ/062+ieKo1
Gs9K2h1vCCA/wtLPqXAG8AOXi3jy0TchH+RNlj+SKFTCVMowHGiejjIRRIKvkD28
EEbAaxJCrekbih2kH2UMF8ZCaIvqY5v7Rf56JZYSfbgTZH2PpyWF/1qUpuP3sjsS
z3kyuUr2L3aQlbcUisqWB0JDshA6X0ctOKjJFibHpCjvymVpe8ksHKN6nUQd1hAU
bhGlLNhLTCrovip0u7kmzaeAPz/EwDA+AwkG+kVM6orT7WEZCpVP8mVAtaI3Iy+r
ElxtrP4CX6Yeu3ZOiX62AdYA42nuLNvzyO9Owb/PgyDg3qdsKhe7qKK4NTqJ6c7P
ggnn2hvtilsv71sB0Nm1Hu2AM8WlEaR2nFQqo6v8TF4tObjCF6KtSA5VK0MtGCEn
DU5fr3uGNeSUwo8WawPu+hTwUv+rZOGOll1hdV+jB5dhhPZcaXviprxEaO3TqfMB
e9vPpJs9tNUE70b34f9slHtmPHKaxxVJusC0Q7OnBb/5gDTplXjcfrYwa/Vwehr/
9suveGjPsgUjtYREyYKJ20XVHx49HIpCn3tr85RWnvLg3RKAcelEDIRQlHFoIyWY
m6RCF4Y3exJqdMEW72i2VWrZC1QcXH00gg8GLkp2G84BAYzw8T5iTao19vfs570y
ccMRgIDx5YHDzPQTPjFNaxjlCrRDmLZLaOUb6edAlPS40VJzG8X/bDFRdTRoTHVS
stpR5DfC19jdA+Prwprq05O0rjOQKVI+/AgWPEmQM2YIzfSBvDU0BAZmuTXpMKll
sjS848mc+u9GoYSCr6Iy966aimy8G3tvT+1QhP0uaTtlhAq4XrWu1rI+FT98hYYr
w8QekOcifjD5xbR7e1WujQv57UPfAKSI0OWnYBBPqqyovbLUezO4kNHgYRyVO+wM
GJ0VC5ZwR4SK1Np1q/2kwSV2qAKoP6d9urWiD3u1BwWh4ArotujRJ+3GEqVjQ8a3
XpvYhs1oz08k48RtRWfzfL2WIfmQCi7gYT8KixkGvs+K52za5ePd0VBCjkq1Qf3S
qfsgeTxx2ptSkVkQ7Hl/giKunw9bXrt8J0/lZ0n5bCLFuD7UF8Dp0/4l0VJMk8ba
H0VPcuayHFclWC1MN1tdTohW6VLLDYRwYhM539i4SDX/Te6TXt7uTCn7AamYIggC
R5CqYT9eLIcuE+GerUa0E1f6/yCdOkpB/KF4y5YxvHd6G7dH7jxz8Xmgcxg5m770
HtblYmKTwfYhE3K+t2YD1iyH9rflNSYFyvcLLR07OatHwO3AfDK0Ca0FEW/tD/CF
xdtZSwa2rZTYyz9UBZ2RGcwuTIgAUGJIkKCYaa3SPkXwu/+xrY1WG4bLfJYkXCw/
6zB5U4nsTusqzHmBiTo/gy0ecyEpVReHeLcVDxHS9/XHwu4YROmdNViqa9EM5Slg
q55mk2kVBe4leybkHGn3Hqr9GEiv3dnEndIHS9tA+3rViCzQZ1AnE0G+/+Ctu16R
elpbj76/R6NAgQMnDG3wb0E26OlXtU7M6K89Cxy5vJa2snau6GWpLKMYgkqjDCSH
UKt7S+d1Y/LAj6C3ftWvartMbl6ZKnKMqxxo5X4fi4XG97fRQp4HkgtQTIlx1VGy
+9nz78s9d43yhSjtT/ZXETjlAFe/yhl5hzdA77F8OLmdYRzUXlYfiJLHGByr6DkQ
dzC4vUmUr/BUG8h72KZi1ieIZzf6Q+D8lo1RwRrRQ8rb30Qze5mrOhlHJaQrnt5A
ykJCB9lGVAQZO0Xz+EwQmvL5FRH7n9WTXvbeAwna+Jd/tpjmlNBxg5BhMcI1TGJZ
DDBGYW51r/uXaBJfVP3EZKXDkm8dEdz45DCgRIsCBu1dmNjyZ15B/dlllPjUDgYh
rB6CatQKGyt7MeTVub/PFRflVP3/FPkLc2+nH11APa5EhPPVEc9CElsBUoOr/YbD
cjxFBXEC1rP4C7pKWWhSG0DHkhNkExVW66mCMhVF/7z/iTBpsdH9TQprwI9tHZUC
/BLo506xMNVIZV4MeCd7qnfP4Rig+3qFvqljUaaJM9yKcd8HqaulpVRPMX2TqBk1
w9tEGCeVti6xe+BiLPGb1t5R0gMBiUDbk8NkgGI8C+W6I/2wO6uzPQGUCoK9VHWG
5RcURiIIZDSvjsbibTj//li9SIk6449Dcc+yFmGy9zUkbDjQrYarapWH6FYaG42h
CZFDQLkt9k7zK+euN7z1f23METOLvXThA0CmX9+Hhj40OYb5d5eU/o2K0zubXQDB
JQwiKPLUFB8/jklGIUIbc/sxQx4Xx2xxU5b2mQGTC5UqsgT6FpmD3PF8pcyjdldi
Bd5t3yOI3yyCF5evgq10bu2nlZuQBgyRM6noFVDxaNaMKGto8L0lNcpjzXozmGOO
3s6CX3qv9lgnB3rXYCTSQ/Z4S++GbD4T4nsRxsl5wTyR5xdJBo+013xq0eYRfUDg
qZ7mndfCnWe2pFkmrvPx4fv7ezsb8qtVvGPgYsCSOX6YE7M13bhwHtWBm+QKjE7b
+gpokF3+W/1FhkZTlC3hKEa5ZGLDsZ4nylDkf2pKbrE6Kq1e0ZBU/XYLRnJSRAXy
iMSVB/ocwLSzBTphUXDoGSdl5BUJK8mG4E25IzKgfWYuF8KsR4NDEqqlq4EhxIyA
ph+TPzEbyYogJ4mc2Fi5N0JJ7xSKIinCzy3W2I8ci5fbN/FNMTsLPSRbefMieEeG
/twq47EhgWJgWta0IS1Da+50vKgfyFwh4M+c2HT3ZqTijEzWwDA+F1owxQLf2Eml
V7FCNwpEjXF286rERjCPmv6KsqWxnN6bUUB21U7XZDK0uJKAdgu+cueGE/oevbCN
3+CfRrT8ZIsgfseEmAHrsgrLeJkt2VNdQYc5AiX6HM+bYhH8mPPVBzRrzAHzfTHU
P/L+9+ihij4tKvFheKvYZZiPwvNQoGxqrr1p8bfQAC+D2Sgm1ooENuquW/J3xHab
rNj5axFqTKh23OQ9s+nDAQAIUikUQs3bDY/0Me1cdWVa3K+WNDihmWHhxaC0Zcg1
q+XzAXj+WCXHLENEMmYdU+EMpIAXYPsM+2N8H5JXioSuV/D2aJ/CzwZrjbUGs7GL
seB4HMCCpe/GeLF8tRmoQ+mXWZUQW/FqATAjmw9vlU1FvYJtjmtNSczay9b5EG7S
HE76pwvlhxX5IRFMf08MM9oE/Mp69EkqxnRdte9FuwoJv5vjedepzK/COtGVy0An
Qgsy2q3L/76Q+KOaOHZ0qWUtD3yUrA8UurN/UhCUE4BPn6UEKU+roh1AozrTELiZ
LT278LYj14yHYys8tayVtl/puqYWTsXOvUHqhth8naVQ3ikQh3kOYFflV2kYvSTi
fZZat6+gnuMa/aAna0Rq0gxSG8uAqu27dZddKUs0XkFpkncDlhiTWqzvgLxCK5Zz
xBSz9AZS9nMaj+Y01ivBfoOydMJ+rWbK9YEWCtvx0p43mP7cKnD7AGkaaRULpVVB
EdMkSrBhGj1gMpoei2dEd8WywOXHtqhuhkJ8a2vLQEPhk1LatmcinTXBNR58CUK2
VksEYAPL5Aoq4vaPuD+JsWdb3VDR/JwP3iyhwN9uyfWAwycvWLw3PN4ukttGgs5E
Xpnz+6bz782j7tvEV5BXTFRSEO7yF60/6Qid5UbZuAgnADYxKFVP/tFm/yqLKKUc
tJQ1RCcxVMZ71XbVrDnXFPP2CpOwvwVihPq1f3Kp0nqUVACN2tEiwRgIjMi4Heob
M+gKWP+v4ECkvpoRzq7y+/MYsAtg/+zQEXNBEKw00ifR9kR+KQppGSk9TyivtuTt
AO6nUBrY8lj/CqPaUFP7AQQ4CU+KgXjRm8eV2JsXdcStxIdkMSk8LAO719x4dli6
1NBig8LfSFKSkBJ4tiTnEmX6p32Xp8j+CaA1BGmaLYsbilR5WW/YxCRaW4/EiNLs
3oTiQ0+PN1Y9Q2BxxRtSH4kDCjxn6OIBBcwScVmCojc5jQ+zMwxt+ZULcjuBe/TZ
OxvQaLR6+h3MEXpSo99XN0akTZkTiZZDFwvD0U00nu7digmzOvTPVe5BAeoGQDQX
QJFS5PZUHlX9z98yGy6NnzLJ6wyo1Knv8mo/uF7jpNSUY3QcScg1D6Zr5orlwZKf
GnbDkB/kIWMJfuqqup9zL69QQVjV+XVPMPFCBRcq8K8AhaTatVm35Qmc0j89ZK6Y
rLGQPrVyi2GRypRn6yTPayaEYFUm48zO0RlbglnbAh7aXQTsOxSRLe35N6S24241
x/QzXA0ZJUZi4Y8TebhRE6mR/L0IsS+jRA5LCK0v+Ux53eBmb7p/khRWpLFyj/4n
UdGv8kFYTkdLLO4u8BEBOBGvL1dMJG3iXnAkviMZgB33hLJ5wPDXRBBS4JNjm52F
EByOWiOnjV1phmziKbOz6i9eyCJ6ofQnnEaNijjZuGgv7RY5yizUSNteOSs09zHr
yJj+v/b4zdybUxoD1NsCG7TlpLZIQHUlja50vLlAJ1PCLg7YzzJN0t5AyOaulwJI
AQYjaaIKlaP1Os7GeB1JsUZOC+RfCTurHiLVqJXBZFylSxzu/3iyXXN4Pk46nVV5
AngFHuK4U1PVcT6eCsbDAKGQKwGk8X/iSFuwFCn3cP7cUvoBFVVkONfLlGXv2l8O
ejeMzJm4T8MstLIzHNnGV3eYfpfo69i+UEIrEv5eI8oq535KffWo/bYQqgS6gtSM
GPV7WCs8/UeVoO5+nba942Bx5Vhi+HJdj/NZNPCqfIP2ckWVW3junJZ301tfIrNu
7+A1cMjnOYnT29ftalB0Yc6Ts8q967edyIPFYE6rupIqXONW3v1Xdr7pMl+zJtpi
5W+vzmPp/N2gy8+/SfCwZpiKiPMVlHN+xmqbcOrU935Y5KpHTFkvIJCDuGAOtzAP
orgOPD7zH5wS6zOIMaW1o8ftx8ayd+BlSrqhmmkFy/qWRaLRDf47l+HZ8S53yoRI
a7oCmgDZEhc9grIhSVceXcTiU+bqHVarfE3X6a6EmYF4GLmvHaj/xih9/wbjVdIV
KveW6677YHmy8uRSMYjst8MM2jksX7ok0v07u2wvcMEOOEKQo16SJvMSedzKd7OI
mcJR4gyjBGwaleb9QTrtd8l+TlMSOs3/gqcLY0+ELxxtRHQFuQVQsi6W02RF39dj
lLwiZbwbdfxMEJgUi3hOU4uycvPfqEzZdhdypiYV9qwWD5EDHXJEt+Ygn0+oakGM
wy6wbTX63bBFAJLy7ewnNrCftxOcF7Lk6bwd5A9X7xrZMowtcMF/MnuFV9LJ/uV6
OylOaixwC5zrUThLCKlm2FDr0MeDHlR5ejvqm61JM84Oqup9QFJY4lqn6VSHtJ+H
p6cukEWJEfRzCshx25uNScJ/WZQckxNpOowd5nOADnFgCbvJwlK7Wl91hxvs/ocI
xq/+TakI5OvIu7DMSFsGjsHn2tiRNvwCvwKKX8tCNz0+IQhHIcJxv+bUm4suV92V
D3h/W+AL0i9Pk2n0U4L5R5AJytl5uNzYf0ccbMJsJCJBw3cNkpuHuWmq1/mzY4CA
WoGL15UggD3nhK2ZSPX2lXVoBouDMLevLc/FUk/hbCUB6pp3dfsrZEe5pbuVFWkY
8M46OJqDhGXEnj3qtX4TZC28I9ST5uKW4+nUiEmERT4xHKJSdYCHNDhYQdc/9FWj
VtVpQ0TeO1AaKsP8D1/TI7Xf+v/gW/OAuhwMClmqE+6w1T/rCaM2Cz7K4+cjxPAV
Pfq8b1ZsYLoe8JlaBNLbbY0aHBEEDMoRTWi5nX1QymX/E5woEsmXi4Xb5qnkrZVX
XJeELqAqRdsXZVYyCGIEK6AanXaEkMnemrMAhwIZsqAR8IgnDE1sEe8+Ej+tvuPZ
7mrgF+94Y/IrcPiKZOVTvKjHuwsiLV5vVlpafQRXKbd5DaJfbGRGNwBVzR6E+ypg
N7n5Q2zE8hBa3aaURhsfeW60otQiangjlnOJL1nLlNq8sJEjsLr1c0Ifd8LL5ayD
gyj+cf9uyBUvmZGbVG253mE+E5eQC0/rqDkBPjB12FEv9mmpIyQbBmzKIDizmbrs
BJ4RzalqJsy5yGESRkO8SkKbp4RPzAYOaos+C0jmltOomNDFxZyYTA2UtA6GFUE1
Znmsh6tZb+1jpKd4wprIJWXQHnRRlm9C9h3yCv2Zy6cv5ZO8lWwyK4JgL4LLxxOK
6G1N7IlXfKHlF434wQk/rxwDQBipVemm/f/VfK0GxgmhX4pYpTVewKeY/SbT3KQB
EyoWJPIFVeHN3bLoXdo7jg/QSA0yiVXYQZqjLp1+LszdQfEzDeoIVCfsPjsorA6k
pHBFS6DB1d0o/aAxBh1lSoxBr7GsvXMhtdwIPhfL7sNjrCWURJM0TRnLnRMJVuuf
iMj+lgSxX/1EYQDobvhBLVhiRJZfkQkHzg+5gtGuae32VBMcWYzv26LsVvK6CjQj
PdK5kKn8nSZf3kXNSpbxzqVS8vyul/ivV2wS9wXzRWjmnlHCRNL6j+YcdaTvxHls
a4uazrPlSjWZqqwEwIHLdVj2rj0j1aIkat5sxR/nzdXsrNEtGgWrDNsLo0CzO1jM
ZAG11In+Kyh9grBl4Q6gb7aNErgteidHQNhBh3u4Xp7kApPldTdDDV/V1UrXG/vi
aSjg9Ebo76TaWx3NZSU7C5WeFpbRSIniMuey45z42RKP3H/UfeouZJxOia1b02cq
ZmP8EBIHHS8d1Of3ouHYurdUGYk17Qaif73mKvw/kCC0QgzJfe5adwu6lOPw16Z1
Wr4LJEJnD6bWuTSJaSCrOe147tiqTq9CjOXaG1nW+Aax2NBOldm0dDpjxrbbyA70
/XuQe8Zxx1IiThvNwmiZsBfbal8ao4QcxzmSiXfSPMLFR8wDUwHCTZtN4FHHPVXD
KLgS3mVjuqeQ65Smgz5oqrpNkH5m2w27ZLmbUhuCcwPOTxpWwP8BRoAMeGqgyn0f
14Eez22Ni4ZHn0TAqQAEajTUo/Bpk/pApIL7pWBKioXE5/mAxAE9565oDHvDdwWF
lxqK7RJalYWSh7onBMOd+16O9rT4vkbtIAN8HZLTjt8HAfCxsWxrUrDHutdjIqbh
70v4MP5ehJPwq0lPERAFUfyoEDs2BdaOflS/Qd5LeyS25Q92ZjcF3HOUW/J5qrby
RWg+rdB29fGjMPmj/Nw+zS5EuxY6UH95/V8++gCIcjd5nky0NGjdOjZFGdgvuH8w
hheynIEslZwzwMSYKohSs8Mb5beNsy7/BQM9+WP8LzNaL7ttzYk1Ni9NzhrO96oX
GhwQ8y1+mhr9RQC05jIBZRTsgGmCn3YzkjmAnZoympZYpmxg2Ozeie0pcxIGGbLE
UIAtWjrOpEUs7VCc50c6ZwwCoGnWfFUrptEroa3lYQSz3ubte10AVbiHsoh3V2pQ
cIqgZoL/XfwauM4kvGYCxzsBRFTStUS42ldhE3yMbbS+5yQzmgLpg52LTlah8lcS
YPtUmMqkZSJY6w0oIrKgEK++13cLZ19e5F0BG71za4Xo/hLXiuW1NBlknjQXLHXv
6LXiNKb/J7toHP5tTQFU0yZVivE4+JFKzgBU93sjYr85OroQ4RQky60QgYqp9oUF
+qJOWrvRNk3PqR0/C7gFmpiEO7o2gdzSKWumh0rjft56wagPQjz7WS0wKoFx20g/
KYmNbC90wzDSEoh4ImGM6euzEQzEreozcFEozmlP1eNES/wZkyWbf0bxbTnmAg9d
tN9NCBUXQ/UTiXnmk5HveQvR6Uoe4M0BE5mlOSkGsj0l0lNAMwwS3bjJRhR0LG/b
Yf6Wjv/51emKGJEta5eJzWjt485OqSZWhGkHHLeixGhUSbKbkS3v6SAue62V8f35
vwt+kk2JNl1YKm6wlSPNE5TsiTszmg9hdifzCxTjjABbdel/OcrB7tAWXttvaqmr
Ay7e/q6UdjyErqmNbop9Hw3EyN4MKXj/0vLMLvRUYIl/zb/DG1U83lryNjB7Z6x1
oiBc7j9rNG0ZEWbN7RqwVWPEOjGRfWpShfMVfBtrcbO0v1kP7Q/CY0avL1wl/h4o
qbCoBtmU70sJD+550KKC+J8fkKIm/+3kpo98qyuMjci11r4pbLZ6Ti69x079BHe5
V/qa9AyOxMy7+VbiLTbvowYAgCrSzxSnBnZThIzwKR/BGZr1KFmpjGNhz3U9m/Af
WeJl7NudHxdv6eLmCGRGXwgNUFYtRa1h4Yje0aS0YG9mbDxod2x70+P7aAN3uQBN
I1WKjVKt0mKv8sYXEOWRIc1nnHH6ItQ658fVRZrdgcrLhVTMSuC8xNatQ8+rLbRa
MTGi/ipZtjBshhGwVKwV1iKDSRgDyWNXFRUArVC0HhZb8PGu14f+BaL9/4S3O/G5
0cNRcO0aqw2PwlfmYyk41x8Hk8JF6iWoztpKWiOSzx56F4i0YQDoNadreZyynfDN
NZPbgOQFeTgGJYvw10vcbJXTL3WXVsBkDOjsOjGs1mW4vRZu7kZKN4wf6GLnEQYE
txX4taeV0ZDo/tqugOD/V8NH78JWg6C/shgx4W/4fXcIYVjiIGWsrDfCz3O2CS92
di4UUFuH2Oq80S99pVifsc2fn+k7fzP8yPV7zGE9E4ZNOxBy0BAQnSdJr4X9X0yJ
nR3QhBCANRybxG4IypPpNva4Of4cfo54zSdDur8qBxmrLSVlIuFJJpogBxzHMr8S
CMQ39bFEqf4PTC4NCtqDWuvWaSSp1icu/aumyeq29U0rnj2sDDWPvPsWR9i57nxP
RTMoEPFaoELUSHWdIGOwOyqLoWdaXjfDWig1un7vP5hUkiknvz5IGQzq8aF3DaB5
OL+LCe94iwUtOgIY7B4pd6U9TCei8RL6MF8dSuapGgCYTXZepYdqfd1mOt8JxkL5
5yR2/LzYhVWk++wOw3ghPn+A3Tojk9+Fquk0s++SsLvGThFIRxOzg8RZzbhueZOQ
cGqIhzss06fFvb6jY3WjO83FSf2ikl5YSbeqJJzUuU3wyae1kbSh66sMBYmN3gPj
ALRCo29ycBDwC3gp1abc9F5aEzvJqDbsmtBtzB4+/z2+rCYWIpDe6mhs3sm7LJKx
C2vi6OcvegOmK8v6qYPMOXb6gTYipqPto+EDO5CgWOPD8cYfHjXrUTNdGD2D4/sF
vKFrDrpoKVljFOmO2pJN9sEE9hDb9u5MoqYu5ITtTaOrvOR8QtyoOdpsFxoP9sUd
Ru5RYZJZfAtYMbN7Zcx81qMg2FxgpvmFgWYxmMdFfBgNr6ullefJGUi5u3g15AiZ
2GzkpkNZdL7hVuir/Tn9C1yr7WLcQqmmipu6l/+BoHDbs1vjQiDw7zf9rmMKToFB
Wojl2MA9xa8QJZzY6b9Tq5iTnW2rnp8b7aFDJfOItEFRjm5ZWkCuxtsqHWMZvXYa
KtkWUe06vlQguNtuoyWVk7ueC4thS/XIq86ayrrzcrRcfwnBisqWmXQYpWUgmDc1
SIcprW6goNb88wSsVnZ0ICRCpPjrYGk326jOeSfKpDiW0Ta0hwWPWZ0tFGf+QUqU
aVA1RpjI/XI/zu7RNiy1k7VSMZ/sVWILtqqQxvNKyji1lgKPRuqqrZsmL2j4cm+V
dVxorPYWvn1nTwc4FnSg3ZqzES8YkBEg5Aht/DRYg7s6uxc0BtqHlabkTkQSP/Tp
ryG46cfEe6F8T3C8RD4mM2IuPMgr5HiZObR1I1AT1+mvrhFFsL+Rnqzni40/p3cW
pKLY49Tj+j20O+MeZJ7Qh+/0LGPPJsl+XAFHXsXFXZp51qTEbyqau2KanRPgLuED
h3LtLvk7AtHp983O5QrQmdl3qq8gcZF2eEdldDQmsPAX4ENPj8fBIzqB3N0H6uZz
MnliG+jo7anP1TueUMRRqmvnOyiwTg0ZpsX6sKhZFmwY+sMomM6KaQ+h78VEvu7X
jHBC97a780aj4bIrIejezuDhUZaqnCOPb1WdKhUKrX9oeEnU6UlQZduY73cRa8rT
bI4e4T3wIqnKhNZ89v6vQVe7utveOOk5rbqr4IPrhtfJLnl/axy2KpUWmS3mr+tZ
HcT10yhnjMUCvriIP8LxKdPEPDCRYfmGJQ+Rz4Ilx6XjKKCgvHQKSCAysERd64UT
IKZSinUwz0INMnGRzbP9lufpYUQUu7LUo0FjXA8+sYEs8OqDMSStQx+rt/w+RNfQ
UHcsCwU9c6O5dLaPGYzALaClqS8JAjxOaIi+N2et1i1qfLPnYLInVB4vxoDu8JM9
X+0jmJ8Glj5OkoxWWHB7CmiEOc1hASi9ViRZrjgQlOZ+bH1CWsXOilDy7mszGGJS
KXn9ER+Gfp2yruVuERvfASt77ksWNQgPKTLEPF414yN7EwzNeUF/NBXLjqh6Zhjq
lhvCe7Vpczx/UNkFukht9eEgj68WmnP+3lGUwOVze+zJOOTGE3s2bnBr27OSxUAd
CHyY466oQEqOl1glDqaV/ea9AdhvRxzjo+eLIWkQrz+e0/91rkcgj9r8bBgr7VPm
/wNWqvMS2l9vexIi9lzFCb9XKTeGFhdIL9wmwB6yZTjyOte2okfR+VWxXaVc3tOf
6Wd5u5gOm9NrezE2fa4n2qeh5vy45RQlVOmKyf/GRAQSIiUM1rVCIe6yZBJDAx9C
p3NYcN2Rm/nYZ7RfV3SP7ZqS3lF7QB+01nmrpGLRjrXDwXs+QUOxhqO55ss0YUtD
FYX02lGcV0MOlirssM2JiPjZw2yEM8wAPtCmGVAQdD8ZuDhSVF+BztZFrMrG7YYg
8HvDQUtD6a6GRoekfKPxeQYesI++ZKuagFW2yrLfKTLJPJXE00MVd5aNwYYwUydl
bxMZKsV2bQeulh5GD1YVgGdlki3Y3ShMiHVqlSA+uCrbCktvs1Xe0Ul5iqSdWMrA
IFFZngNayIIpCLzDIVR6JywWKp1hRBsSXkQYNehKlVkQqwlUSjd/XXXFS/vWPePm
mgP7K5ZgDNS1etmkpd4h1zfeRqfB2qyWLRhL+ExGlOlwtW4R1+q9RxblthW5d0Ft
oz/0Fa1vNgLfQhjbuTLulnxOit8N40DgBJTwZ//8d2Owe+jdw73dnVTXcoyB5nVO
h0vMTFBBZumIJJ9uwIIudZ64v9QlvHSO/fZCXVrzXUO3zrcbOsgHRJjFhfAbaHex
7H0G1mGbkYt0ze93jLHfBXr7jSLqYSzEppibExvQ5j7+cDrrLo1VAaREdwBxA89V
OHOX1jN9LXw9gq7qpLjRiaLYdgOCBlcH+hUxPKlADradJ5PqA50/mcTuwWOpfSps
DcTrpM2MC1UIH7vf8cB9gvHXO1W8r2BfEWAwYIywymUy0hP6GGZb3plZORLXWYfx
xRwGEXY1LcEAve5HSfD0e6wTjkBZOwXzfsixCYK+rATYQuJSbJiu/tSECBIM75b6
Oh0MOi4DbVs/vuHTekgqVdoYg0tdWPP2AluT5aLUGSsv/UVmlCewO+JH2daj0mJx
+sp6ATW0mxMcuwyRDFPwsli5Pr8a+93Ld557lkPTM5udZPTH7P55USBT+lMgRZZz
P90K/UKdSCRl2FIG9D1LUyH8fXRgwD8E5jkq/NCPuVuuOiBPxW90lpNVGHpN+OXQ
R0oPLsTYTRzXWBOkgKiB9ScBXhCfu28MTXr4OK6RBF24aPBJzk2dipedBJm+/Mzm
4LWPDy+e2KOB4KsjoSCSmHdT6o3WOALy040S8BwTJtTUF7CxHfdi5T0mdDdtJJsU
lldruBI6kicXPRoGvZWC24MSlv1Wa8ht+1aRu4zLu6Z5kKJEC2TgR/8/iQGZevNV
n3vPMmgAUd3y+eM+gzIdk7atBw2EdfP2B/eBdEL1aF7g6FFQSwlu+TVpZTBSJlQY
80Q24OAgvXTxe1wQ3In420Akx8lglbI9hBHjWr5tMCTZ/OKAsHOcwb6P4vhmyjIb
nIjDrHI8QzpuLuYwHDtGiDHT91uHSH3S8iXTL3Krm4cqvC2H5SwOr1BrRHwfQLfY
W6p3FqxR4yPxqHRdhsMGCA1IzbxeqQJbMKNqWnFDeHrHcwDRY8ncsWaHMiPiH2pz
wl48gTbPwvlNsc7/QgnICvhJSuBd8jirrIE2BaXRxTIXyczB7opoMBrk2eH962uW
C4JSNoqFVHNSmhIeKcxaA3zFP7KsjXEYe6YSvDcd5ak4bTfrTOYpjfC8zR5byGI0
v6qwbJmV47wC41gD87AK7qX+ySGcyzyNg1haToU4M2N9iiLnsw2C1JKxZX0lSKrs
ggal2WfglkKtBZVlhug4pZAnBGDxHr9fkS75mNrh9PBKwBw1C5DaD5lDbxBDi5L/
x3ryMJKarycu/3vq21Dgr1FoXFepsErJuwRBg0asOdI5X0EI7AVyugBpadftZYRg
UiWhpjY92zyznx0dvBHuhik7IEHGqD7exG0ZFggE3q7TxgDPsRfQ1F3RI3W79ICg
eJJxBXPHW5fsx1utreqvqNB6nRWuXJJcDQX9RTrv5xFicdH/amaLM3ie+SV/4ZoQ
tipYJrwezHyyNG+2zbfBJqMZOizC7FwSuY68PDLMWpu9Eicz0O7vUY2XWUgrXySf
YwhAbFQpPjiKKnlnmjskIs4blG57n3xdg4qNAkSbhWZyrKhp2hs6m4JLfLnqRqRK
VTvD6CUks9G7oiiBYl0mcc3+/89Nu4U0WN+mt622uIKhKpujOP3ZzwDM6rUh5Z4h
7TU2y8WuKXTGRY8EM/9Wsov8m0a+SEMkL65ewCwNHu01I2QQI7HbgQ6+l1kbKBqI
f7UZqYzOhQfbY2oeHGAFX0vjFK1/gwj2dnCf4o7H6h63+Kg0zRCsrvJhfTN6WfLv
nmgjb560bDVodeGpJkBiOFDl10R2f4CPAA4o64p5bWQUh4dS/6XGmncjkU9kNZHy
Afvaoasg64sZzHl6TXm+3a15zSF+Q7Sv/m0X2KTUCDeczvruv5TpwnLOyhpId+1G
Z4ylPgr1qHUlwcY3QyPRU+L1FSpfFBjUtfDXSwLuuIuKIHuD2lWOTy+H6krQfVdD
QPYpBchULqnj7ZwTGqWXJ+bqD0z+GLa2W93q3czceFQuamBJYhO9U3OxlT8ealpn
pzfB94G8Bq+XmwVZxWbxrOki7nha8H2D0/zWJ9AL52m7goGPscRlEE7AtolgKfTE
OfK03erCDDMgHxGn6OF6O6c5eXikQe5dyUPU8lDi5c7e11t0m0I8iHeadACAbqac
+KjajSkWrsXysO5gJ1PIQSajhO1kIv8lwnIAas3jo7Qq0msd4mwOeQHujuqFhemf
Lbo6Ep97vOY5c8dBFtvRFUWoOxvnWLlbpeknpMpXQCF0Z2hi5SAHjmx3VA6aycxx
3Pyi4mY6VkhUBVBiZFCt9HSKlPU0Tt3sdieX+xb4Mp8t3Ab9bbcRMDMgTBHLnKut
cUSZxmb8wYyfnFd8f+xGFXS1HmtLfAm1GYscpNuAex8FBbrhgHQcz9xA9sq8JC4M
Z5XXIzGhGlvAVIdUcnHXZzrLGp1JXfklzmLG4/mQfrd8sc1FkWKgqi+5+9f/LcD3
iyQRevXBLH+xiNeb5qXx+xyxjBVUBrDEo4NPFkWHHYFXAXnWWoqcxoJ8/mkiLItT
jYe7Z7YkkLAUm8IRI6Wd4ppsCl/Hp7UElo22tLfDwquFntVJNcsrL/88qS708+F5
iZPUAr1GQJ/NfFNjwqcYj15/GakK5OTX6LzMbfSon193cxqdXAYsLEDG/Kkkn0Xm
XJ+BF2aU11IOWzH/JopXvnEw9bZsfOS0QeQXTZdxI5z96OmJkAvmSTVZGU33MoSQ
pCq6a8k4tkqY7tRGdUKXZu9jeoT610/iFZcMoHgpTdS/zLSVr5XkdC0znFwRw6kp
ciFNciYY6wtDp/QbdOTKLlLz7l+I4araeG9zjtYZOrszxiYad/pqybnyRX4GSQuH
zWKfGD3nQyyf0cvFd+vxvJN+sbaFouLVRy7WgOzks9ytUkGQFhtpPvEuJgiD4CG0
79B/X+84yBa1aiNqdOkVE9OyfXs1UR11q1Wlr2sXg81k2lyc9zrzxT02qmhFQKKs
psoTGxL2sAOF2Q5qHNwPSc9gQM2+b27UpGg6eHhRJKnjI0fHUQj3BNLpquuAF3Gf
sEjPmfDDFnC0lSA2/7fMwE3YywzPM53cEpgPPxreAPeq/96Dtj8OHyRc4FqdNTM5
8jR5xuqg66i99athYxUx0lIhF5MDsg9+xfSNbPLYxJjLfDy96LaXSVs4l9qdNebN
mjruMIOQNMCS97u+J6LHjI3gxVb+AjP1D7JFgjU0siIoXAuxQ65c7hmTIoIfdAmr
vJlQm6y8MmW6wdqHPkmJUWfpw8DgmTqyr/Pl0A+xsZzPyXE2GwJaIanLiPbYwQ1j
AodqY4Qekn9txL9g6VI64BX64Dy1pbrjG/9aaXrPNXZtb/ccb2Fm/wqS2b9GPWhC
5m5nZmtid9E+iUNh4NSxvkPERNPnD7yLM3mm41bCnHnTMh0eeWwQZYzM0yeuMLIs
V7IE9f5ZoHwwAsa1wjTc30QjP39hTY1GWCrDzM9FilbVkY/FaIm2d+HUIk8l4ddS
PJYUuBTsVe0swq/HKaJLVqdcbjsleDY9ZZgEMDsFmgooTl7O7lu3iM/o/yfqxG8u
GtiqsN2RZUbqZ/OSR0QHIO/iJtib1z5NcH+SpgSUw96JbwIYWSz37bcGTkFTtiPw
hxYIolu0kA6QLbrkPxjdWmHxxnQTqqyNxwA3CCw1y2lvGu6qU2hwdx4Wab3HekVZ
ad/uffGQT0DGxQuY0YZdDCDDg9SpgqBm0H8RTKne65kjYwdyeWj+2L3/PW/01CXy
ZBf9kDHNxsdseUZhjbdZFUqJXhJ4Ex4klKNFTyLyOtJ5cLD8rTyKd58eU5v1Z9jJ
EC5Bx89F3CphPf7qcRYELFjS8a1wGsCdxxVUrdoezVZOg/Piml0fBlj1mMgkXpwg
3a1WRE0URUgTqK6LYET+A4hbCzu0IgEnsjxCfxMD2rkqXXD8GdO+5CZA0MQcVCHH
03+mfDFtMG1LUT2bjMQmBLvLUcQoTT1eIPjHkich+ncjfR7G2YuPpHKIUR8qi1eB
wJHVdjzRaaudZT3qVP6eY+kHJGKxeC5eneFrscYRIgcTR9p3rHBb2TMM2uX+tqcL
8k1Lpcs5a1y3pR5fc1KInPEqHRNv9vcAhlDHXKGwwvh0y+qAQRFLvxcI7+eELZKp
rsjYCCnYscgd4ByPtyHmesJFCK7cQ4jETskzxfeFN0NFDZjmIWPA5p6dDfIoCvQI
ByoBBys77WeGow11JqkTbY4bQX6owp/qiXGSW9hY8m6kZ1x8W+hVH+fv8UgQE+9v
5NCKPMFQkn136cCNlhQB8SkrnCrdoNTUFHD3PC9NAcxNMv/8d1IXxq3EqJ5v8b0R
mCJmepREYknsV9ylor7VfkQP3j9EmFiV8FIqfSajf93WGIjIAvkYe7SJuyZPrJEL
Zu6bxNx8kPamMiZZey+hsvzYaXt/25LQrSYQbhS4OmnEC9J/nxZlmI78ywx+LmHw
z+EwF6NAdrHvCUuqOUIvuKPIeCk7Rz2Un9bCtFYO6u2wtQDABuaXdI6w9dkkHihn
rxYXe2y4QbU2mug+ckOhPC0pqfgppE0AvXeGYAt8b5EKUUL3VK33l2b0AsHwrhhY
sJlzP7ycxzxDgQVHAPBZkXTzgRBKis0tCLjkX8kTEMBIAnUbr3T25yRGX0KF32db
QODfFeeowd2VhUYncGchjLo83C9lX8Zkudem4ElVJf2BOAAxHUwhxtY3Xk1+NVf6
F5vl3tOJfddegGURSfDmdh0v0f+PgbruGJaIY8kh+nZApIP19fF2wo5J3mdEk3sm
NEyNkEABR4gj2FkunnLvcZBrZanN9+kO8K8N4yr5Iy4S12wadac2O+NO0RxcLIjN
hlZ7V0o+3/ICCRnLv71eARbFmWxwSjt5QAP5fVWY+Gzq2vFWDfhNsO+W1E9pW8uk
NprR1WUZokDa1KcsM/9g4psZtkbLUmHtyDdw1PFobNVwAPcTPVfXDh363rcHq7Qt
EtQK/xyiWkfbHfF+fp0tdG1TpB/KwY+BHvXpmjrGgXTwyan4BOx3VsMu6U6i449G
zwGs69dq6IsDw6/d3Yohx+JiFLpu3EOLp4aTOGRQFnBz6mnINtHKc1qPK5v3fz5Z
/bavuTDgkYACJpjuF0S5NazbgLzaTNv4a9L3FckBvo3IMAcUShsNbFItn0nMYvZA
2+clPOoGaa6Y82Atmmc6U5e5jlF+K7Z7REL2uZ6XySKxBY+YlcWSosU19D3ipc+x
r/s+C4kb2lMeGb3dveRZY9ixwxG9T2VSRruEJL5CSO/1pR3sLrgYKwus8qmAxo79
1Zw2ON72H+uBGT8YebACjQRXTUoJgEAvkQxgRaeR+nstZaqoD4RUR/XZZ/uvyPJK
KKbm+BTirIxB8XdV+TCxJfovi6AeLiOJr6v1B5qsnbW/TiWbXq2/pMaq1qVWkErl
fs3XoRU3dyNhGml30sSpzOBM81aKa0o41c1XkWqlJZIWoSDBMO1tAETI4qZZ9Z6X
gTtgInYX8PYrtrlA7r6UOEQljIx/PwCilu+iMgMn4y+oLEkexTU9q/txc5U9xOt0
WUTmuwCGNWGGqTj8N3dHUZylMe7Q0Xt6R4LMY5w7/eojGWol1viW+C3+zuHBmXPq
QafqaWMTl1VD0A0sn4NxoFxXGVG9pxQiXoFP4sVuGD/osZQ4zNXdjX+/U1tFWb9O
7M0OXpGYNXtp/EaZzEWo1zfAm76zBR+hjPeWhr/dIdZ5R/QkO2ZFa4saVh6U410I
BwA0v6BWC6jLjMIaEF7Y1Cpx1314pvn9ny17JO3WbH6wd4CNWQliMy4TY+FX0IFm
5b7VoxE/gGNNa+GtFRcIEigy2K1wpH+xF8N+KSgPZTCdeaj7kuLxAhXQhtDQF07P
yUx8R1CdCjYtMbQ1yH1hgcqg15cVjte7waKSHWgI7LU/Vxd3nV4LPUSBTTmujc4u
f3h7z3MI6GsW/QOnl+3P2ry6x69A0N2tacwX3mT60m0OUZO6bBLxtd2zwhCJaDhv
G1KVpd09emJDtSfY0e98lhQzr/P13HbdDEI0ikuHTfM6DslinsaKsgX5Bju5wcVV
MwwJCwT6kkaRvW4wQPz36vLqqcCllaswtaWXg9kmIYrTGPUhp3pegZR3PRrZQBhX
pGy5mVcm6r/3QgeTeegM2XHEs4yFQTihbREehoqMPgKpBjpSYplHp3wElEUiaLH5
YYkzux/t/B5+wFemXbIPKKVFhYMAfdAfvgBviOiLBDfjrDDMEVdqXRQhylr7R0I9
41R7Sj34fB0aCUxAiXglpdvPe36bQ7xXjh7IPGoKQuz2PXowyRDxRtdWIMMNtALK
fsiU01TIPKEXg5GzfXSO1kIdo7xiBvqYh0tRdYR110bMBgiftzIpSWmR9dWsuQ+R
6TaBei+ibex2NwkRjKF9eqLkZLZ0aTLDqAGS4bOqfhSXt/QNDyibuAHIYssIUmOI
6CeKsgb3gE8szbE/3foR9q9Ek3izvCcJqOXSv8mmBWqOucPI/mbPpg2/G6OW8uMT
NayBF4o3qqd2NeHsWChEvgKgOvnyFa8kB9g51AMbSU2Ovrh7jo2Et7xiS67RU3fP
P9P8om+CAZ4NPNrbCvCOwfX1J7BmgZmQED5RWdCqsQclcftAK/q7FAEris6CN9YL
JrhDnmZBmz8D5GO4P1Rhp/pTMqMKXlwiwxUNz65zNmCGGHy+RekV0xmpGQ+Xcf+m
ARMT7DIpbuzXuj9XDVIbVd0jvnFoXBMgWYYFertHGRHYlrx19ZLqU3ImsXFPvTtv
w1+ZPdaY+sxhDXp7Jov9/chV9+emQVcwpqNolwaUPUIa9EtEdEVuvgeHb5rEy+aA
rvUY9q/AACIv7K78oaZAeX+uFXJ7a5ItLSHGpc+4ZY3Ky76zi0l+z1sqpAFm3UVW
xAQmdO+F3r32XVA5UwU9DAAKIDn6J7ZixMclP1n59qQNV9YJ+9EV6aVnFwhP18d6
1t6cuFT7VUyXsx0JPQ0uL4qoAAY9XAwloPx8zjPMqM9udPc44nspy0L5N+ATyw8Z
VAkrXxFF/ImbSEuqxKD2P08cbDURLwD7jBWSNyzoscZ8W2sOlpQJTJR875nGjHL/
//pragma protect end_data_block
//pragma protect digest_block
swV7IS4+nCCXEGvWB7Myj4rZhrM=
//pragma protect end_digest_block
//pragma protect end_protected
