`ifdef RTL
    `define CYCLE_TIME 40.0
`endif
`ifdef GATE
    `define CYCLE_TIME 40.0
`endif

`include "../00_TESTBED/pseudo_DRAM.v"
`include "../00_TESTBED/pseudo_SD.v"

module PATTERN
`protected
[QU9WUR.MREd7MX9AH/OQO<+G>8QbN_ISAafgR<E>)aVA#cIP>WA,)/a#_OgGG5;
I;(c3d:&+A\,F,2[fL,c[(dIIR)EUb?9H=<e1DJ(;0=.\^K]UL\HVD4]@f0ZD]2B
K/aN/\0e)P<K>7bP@LP=5K#CC#0QZ?I)KNc019L-b5.C+8YK;(YO4YVTYF1H:96Q
8AP49>G4V<>D6U-U31H:2Y[D3AO\.K(VAVOPSg\XGYdJ;(S:)UZgCJV48,VA_CVG
+I4IZ0[M8_V:4AWdJWeV@BG^WeI\J?(GN=>XLbK1T^@+DEbFHC4b;U/UG)Y>,CB3
fO,9#,RECT73b@gb\+^;PPY0O4De^UR^S-LN[6\^a_6N,C,,HT^Pg5J)YP:U8+=8
c_VZ)fO:E#CZK1/E[P8WTO12aYG@@R:(4dS>9R]PITUF-TZ+)c^_H\NcY:LW.b9c
PNBg2^23)CS4(=ObD@fZI.Z:Mgg#UU&CL[]&@=?L&JLN(3>L+26?>\Vf4X\TN2O8
EUc+R#+SF[+b7c[.6^)@BJ@.O05)<Q#7OJI,U2B_S,#\@<gI.(b,8OW[[?<(N#g,
4aC>Q_Wc(^^I0@[da?AbWBaB.^KX]L[]6cVWPT\)52ZA1^_IB]];EZ?=aQRGgKYZ
fb)Qg#V)9dXC)IKW=B@6f&=ZU6-?,6H6KHN-,N&IL6,K&8SH\1dSP.;E7?/fO.C,
P.(UI4>9b(Q_(9a520b;GAf603DJQ4-WZXb#^8ET61.W(DV5SI,b0e4\?VKU]5ZO
&e(5GaKLRdC,[=+_&8B;0OZHaFCW_?#[-.6/KJPE._HQX9FeZ9>=ZcX#FQ(5JbDU
/=d;1BWZ[>fN.T4RFcYFeM+D-FW(<C10_7:V]JE;BAETJ?4&c0)5QaR#eb)][.XE
01(+62M:U\N?IIZ6KJd^061?@KdeJO+9X2=J_I<6d?LQY0<Z._<F[#,cXg1^?Q[R
:bH4gfN&R3NZ0N?MHO0OEC41\#RM(AcZ_b&aQd[)fF;_YLXJDD)J?C.f;gY27]P?
OKN80EQ>:6Lc-XZ\f^;5J96^A/g?33F1&KFU<d7CEOgC+W8N,0L_=L<8A?dC-VS4
]ZV(Y-GV9?F#;.#([]bOdF<.bJ#BYP,2L(MSZF4@EJaIHdOLaJSU@3/^9g43U@XJ
cLAL=<c6DDCb#&L^BgcNET/Z;R6MG-e2G;>eF49ND43Vg0F_2[=dK6FYSWM\OIW(
X4Of?\WQ]D/7ec^UCK;)ab8\?fA8.fY_FJO0e?2RVLbaC65[K1&@dZBU=#eYG+IF
<^;=N:62;a;6K_05SI\.4=-0bZF/\UJK]Nf2BDMa-6+I6/XeVa,VD76Xf94,8:_<
f;\AA4e>CHFM4>4Sa6Y;ESH8:TQS\.?@fPV\9,M,)/:DMPI^JN--Y#4eaG6T8-GW
:Yff;(>[Vc&30^7\1G;4JY)\9#DbD-XNA7,-0&MH+K&^/.&]MODcPD^<.ATM9NWg
aMOYXAGT]S(OaJDV.UK@[aS_:(^Ce45cId/eG^FJ#Y#M\^TgBZ_OXd1BDD/MXIf(
ZRB0f]\EBA\]YZ66LDCBa-7D0>6P0QI+a<3=#,]27+bOcY^a?TYTAg=F[gHW;5U;
_N6XQ=_+>&(WC<.+fK98D:N(.eY&Q=RXI/8dDgVdVJ:-3a=YV[7f7X,Od0cCBB-f
IHP5?[,5bJJU^eIJJS(#L#cUC7=0XG\Y1MZY?b0YX5T,KDg=F<3#ZJ@P:9IQ-[]C
BT5dKR34)8H;W&<d<^dQHLTF1L:I_V4Ug)LP5X]26N&VLfL/ZBE[7X-f;E_^UcbY
+=W.bPY^_Y1IC(:00X1USVFP17dWY&5>a>A_,WE6eDQ)3HafWR(f9\9b\=8aMY_Z
L8c3\MUV8aRX)Da=JbHTLb;>(;F74RgI\bB&f9Af?QFEC0eT432I2E2bLF<R@YH0
EH:7f4<d2>GL0O9&H1X.d0=SSb:BbO[Rg=:^6,<)WgHAMeEL[.?_La#g)fQM_KgR
Y&S\8a]7;(f_Y76H1V2M06.&3_aOfcA0d#];fe//?A(ZS_PDAI2)&,P]C8f1;\GM
Qb,b3H(O-N.;H;R/G-)bEFE<gO>6b_GeKD+6eJgDQH[X?2VX,8/]P:X][8[NHY2L
M0.dU?\]@]3MgcF5TMB58Rb,c)[<4\A5cITD#4g#,4X,X/.L46Tg6RV7RLX2P2IV
c5.Hc64QQ0FFfY;8:Tg6[;OH>M#4.-W5;<ZFJQ>,cI6<BX^fO:2+UH<6aNX87NJ6
1UBNYb3^56bBdG,@V<>@[86.<aO,8bUd?6ZYgG5<[Zd_NLdYH3C^c9cPFU[XI>SK
JBdJX&V>>)69.2TS#I3.K(L1gR<cZdKbZ1XYT+K1/3cF/I[>5B@bL#JX>CTI__>8
e_Q(\Cc:7F+59,D_93]NI?NNP^#_1<.PH./3&SY6J/97a5VO4)dOe63=OPVR79-f
;AFaE93<+?MX+Q,dZE@feN;GdK5GSZC,AgIOZH75@fd.:WDGMa?c)GON8Z+=8gca
AQU;O:LBY5-)7:DMI-eRC9T)Tdg\4dfAIE1V[[I3J3+3K>43bB?]YCH__;RR<\P&
+61ff]RWMRB]6fBT,(,<aIB?2Q^=Ae@:5<A<O3UMgZdB]bU(.Q0(OD&UAD1520WM
[Ke=6CR8C7d@FTET(2,0JeI^KRd[F#ZS=1af.<=U=E=g;VGd+b5UM.beYM/7D[_H
CWEF4(L=.9]7XXd,,SQ=\@WQSI8-_8R9<VMV,2D1]J3OS7Q.c5E.=\e/SHdCN?[;
U@,eP\+WV<:a,WKK:[H>eKDXKTg&gRZ(XGO7g,f9aOVGfG,IRA05@EP;#S@<>5_R
.fYf7AWTKW;]Zf_=D&4O[>OZ7_X,RcgUb)AJI]3VZUc=PTd?DabT/0eF+R66)JTO
BSdRd9bF>b4(Y^PDWe.I^]cT6?T<TEbaPY5d&__BPS@_LBB#^?<R69:(1C>>d^H=
D-6+0fFGBP)-cWE(T/aPM)U#gF:ZR0CL)9B(SU?aZNCTeV@6H]+KC[Q>(+7#.d1;
6WN?J:EaGFG94Z6?,eQ?dSaMCGagg\EBg-9FUTE1.[LLIOe-gLO9;d<S4b&\[Q#8
V9:g=2Q;?cI3@:D7617O83(RY+S8[DD^+N[fC8.@;/X7Z-L2Z++-DWSST,,K<;/D
WL;B\)]]Gb<;:?XS99]L#7S\9.4eVMQ2J-H#\JP=&I,5IPKFS_W+4d?L]))@7:T)
a&c2P0(M<fSAT83J]4<<0UQ>9Sd-/Dg,a7aKc@G4/fRO]E8AeX9XGMa?4W17LQXQ
]^=DgUDR;6@W@QbH0E6e[4I[G14(UG.WN=,fM(VgNF\DR9=BY1/TEI0.gc<EO=dP
W,fe&\TKg9Y,K3WbEQ&H,49P.-5D\@F4<FeKSd[D1KY825/H&_G6SD_5?JM:<Q;(
&H\FS]-)-&:P+49[VJU<>&(TBK?56L14fEQ6@Je?G=3fD7<_FXC5bG;?@#N4.&KL
TH6+Dd)Q>GT+^Ha;HPZMQX730+U&F1;+\\IA)KY];I8-9<Xa\4[2:[TMG@Y&6Ec9
NZ07VbX44=<?LVaDE.R1D)CV<9KdL6)C.:ETB1[F)ECIRDGN>:[R[dFg<O;W6-[<
TX2Yd8VY.7H1?A(&>@/;,GGb:cA[Ig\C:<&@4\4V2,K?)B5.&TNgD?Y908+9[^Z)
;4<.I3#dNd0T.W=bK2ZY@edT\)Og0B3(0^<N:X;Tb9+(beH22><F^:X1+GaP5@U5
5ZP@,N:=\fL_E##BJ.?HOBO#BL>M>b]A&3=<MZfLC5\(#,g/2@#GY+W0.;F=<c:U
2<?X+G.:E(]35LR/eNPZF?)ZDM?DUIBU4=a())&g-e&7(@@3a8]U4Na,[U6[fU_H
CV-0\S(U,8#dQ3OG4D-M5EMeK.ba.^K3K07f)MfJOUOH6IF7XRg\+#HOK5\dD@8O
28b3TLgU8MfdC+84Jc<(MCW]??CHXU+KNG9cU;RMHN#4UaK&#+89E(G9d5X_Ia#L
[+L84YcCU0Y;Oa?\dR3:H64CV208\V/7X=b[8L(ZOW6,8ZXP/^R[2M>,_OSL@E+Z
DHC<QgG38)&c4\3GHb-G4QA;Dd[0R+YZ2S-L?XEE-[>33&2HV])NV.0CHc9STSZL
^CO52;cZV6(/.+XUe9]N#D8NIb?,SG?@WSg;ROgJd/:UK&OGf93/LJ7#c^)?^K&U
R_\^F8OWZ4/=8_J1F5DX,e1;5A5gJ2[##5):^^a9LWMMV]gH#8O#&S?GH1D-G^N7
gc8H,4FUTG0(G/^VODCa7#g->GYM.C]0I(=\O@Q+[eD+JQSfW206N>4D0E:CH_](
GOF;#@3AS#c7P4a]7e&ERcQWB#VARIC\N8.[Y70B/R;&S<X[,&W:H]UZY(KL7Se\
Ya?6:J>AN,/E==O(H?45c;.&#1W&2/bIX4JaI\+[aUYM>?6WWIMM2YR;0<e/MX<4
KH8].VPK#ZbUZV[F=b<dCU7f8UM?GgOG6/>g_EHF;e^]1:YUFJ+Pb/bP[,ad[R/.
EK@0UZ,Y?Ndb+@@OO:4L,C+N&(9Rf.KPA/R2>ZWa(V5=>IJZ.0B5_,&BC]FJUeG+
]8fJ[f<5/3_L@5I/0.+@&0dX[AV][)K]32Q0/3-:RBA^Q-_eLfEgKP7(TB>;f\@I
,a=C8NP90-e2g\gYE4:Z)CBH8349SKJFLg>4]3C-+f-K#3MOV5FXQUT9+9&G-V([
Ga&fGg/6^<Wa+>O1XaZ8&be@6.eIg:1c(6F#-<Q@D&fB2S,_ZHAR8A#\_1_TNG&1
EN8Rb,WE9+^8Q-cc<6&JfZMVN]fbO)>FA\<;09@8U<K&E0PI.9[cN]G09)BDWa_8
184BZ64N&.J2f#[FcF4U[&29I5>/(9I]VI?bc?Oa#W/:A;EWa)6?]fU?E\NADKbH
9/8Y/81IV.0HI+.K?d)W0Xc2H+;OLKD9=G_#V#UAB=&aSA[TWXc:a_9BbP[?:Gb,
@]/[N(GXc6YV_J4O9WEIU5FJ#BZ4W#5d?+V;eUF3=e63):-#;A;]HO2/FX8SgWe&
/d#V2/K\c1@UO63QLUN<^YNX6YDE^5+.)70<CY<c?Rd44a\QB0ZG^\91D:#=0T;G
/CS#PWYPe<&T3QNB8.2YBNGQ&+28g8@)MS2,B=4\<.5:IYQSQ@_gV8Z/G]T/06g-
V,+f1Y,)P@Y@22.R/ef2@#^0;:7^30^VT?e6(O&LQ_(\OEd]6-S&;-7)RVZT\Sa\
^PF#+[APWJGD#):0AeNf[&C>G45T6&@)RcY/f5ZTL.TZ/R_R7SR;>J[+@<0X:^_X
<WG;5R>:ELN(CV-D4[9.89SS)OF(R7+L7A.H=?XI+7J@DdB@R8.-X#BZF-(V9b]J
7Ab0O4@FUb1;M4AXF4H?K5>+/<3C4L5D:V0^J(B,#[LCHeDe9&Y)^O_#fa)6&Kcf
[HJJO4D(4^1D9J6>2&B0<)].=[VO.K1MJ@1Wd957U[Y+^KMD=WRLc66Od7FMVSPM
()M?0WbVCA3=_H<VHK@X+NL32&:9JaV7eI(YBLg\?_@He&NGJAXY;EZ>cPJNT_3f
e&Z3/]HB]K3[BBSWQb\/>48QUD^#\C6Z9TbdH>e?BJU6TUM/;HeIKbgbH\:G3g=F
]&_\dMU\JM1]<+20R:C15Sa6ISb8LKf)Q)Ad=a@L5>LUR0)YBZC\?+E=W5g97G?,
-ZaV5KLe\#QeCd/B:_;/<E>]\5/MK)X4e=9@]Y[F,]B[)H&e\94_J)VM1^J8FV.f
Ig15127gXN;6Q570PR=HLF8DHTG=UW),c.-g@<055Rc5DW<a2WJKB&P;3(#c_K@Y
IRS<:DG&IUZOYI-8X:@.WJ[L;,c0D=#e[TO9V=2PW/f6YZSW/5cDM#gNE8624/7>
29RHB?E@CLNCWQQOZS>N@)_a6ODX9aFIHWdc?/;VMI\S/-6I1aHbcF0(&-3//H&K
ZO<2&[aLELZ0bNa:[/K+QBAWgW=K2MSKbgH\dT.\U1eG9b2F9WWg/;@R/3Ne<@,2
;52WRGUcACXM1:WB#PX_P.U&YHIg<K^e6272Hda;ba;eG,8T3LS#dX^^SJ^e+B;f
17IbS#8_AfI.3:+5W2ggC]fGER^G\07@1@OS??C8caGS/<ad;.RX4WYJ[K:NO:&+
R)93GLgCNg1KdZMC_))?L_^MfXMN?[QeaEf0M1FTX/Z,<B0:^:XVb/g+WY<R9ILJ
_][a2=f-T][2O88SM/R+V_JVc8]df:7d8<eR[AO2J.L>eYHXg-2TcYOVN1FL1NE@
^AS,6M5D<HR5Z24]YE[).Ca5g-8:1NYVUDgBMHBL@PPP>+[OfY;Og]4b()3DN^\J
Y/WJcIe)g-/?XY<@#;29\eJ[V=N[VDH^K]74^G#7Oe0ENKL-LW_CfC4K9>YXEf?S
S(=(Cc[HJODM&WBHa):#4Z\#53O9GH.f8;=W#27NN[:]=e;ERM>S28VN^)&.>FaF
=aP2I;8=;g;W)^M7ReJ7JXI8<GA;W2\EbeWOL^V.A:b+#^8DQ3_Y5M4DgNRHPPN@
7bHOcd:.d/_F]RG<cK:UBT6/U\B.c2=XILDOTM9a>IdKQ+cc8+@PQ\,<bf\(e?-@
DUJSfS54VF+B/fcJJ=EH#2de1+A-]c)fe7KAVeX?3ZeMGeI(=0G,]26b9]R6<K/,
:6e(DX/eBTED8PY<?a_\>>_BQ4WFf:&LHA8.THWE;@CB00a.ge8Nc=]]SUVMK7\A
Q]@f[_E,-Y&d-6M?6JX5KSZXGXcWI\-(9C(CU<c/,C=\[ScCcS>gZ@>Od/<A3>7N
?+J4>],SZDO.1#.=3S4MVE^&\Y0PJ2I5XT#B;R,S88^3IF-67=OEedJ>@DdZF)(+
_VBJ1@/=.TFL>>,>^X?gB<F(]dH=c]-Q8&]FP#bOG<A/I)IM.L8;\H\c09GMX\MB
CR=4:;@#-7AeC4J_gP]89N^&LR1O0W-\:J7fa67963,bU;0fLfW,I;CSI.4SC@44
bNW]L0L3HIAg?CTM4WHbFWUXeKT&DgUb^KE?7ZA;&PW)J>gL9C#RZW6+ZF634E73
\bUgaWIa>)dU^<<BI,d[X)H;YF9YI1:U<[A/Va^-H_Q2VIfOM+CGYgR:M@IA>NU^
CWI+]3cYJ&VT7:H\d:G@B-=U..XLdP.#\;cN:.G5Z3T-,b5g-=ef5@GDE[@SaAg1
F>@X3=?KPU<]ZE&^DM/-P08<b2]gP8SHXc<W&M?VX1TZ1-cLFDPXDZVfE2E=N+)g
bR67@.+0Z+YdR)>KGYBB30R9^J5C3-X\A9b&:).g2A<QZ.ABe4P;72&M>>UIRgeM
C;T,T8KX4<W5,]E-OG]g)c6OT@WfRN5FANIZa_eZ-QHKPCE+/(MSMMD/G9Ce(R&N
fY9I0G]D#4@>gF8T<[.W-;f3I(U(&?-P7ZM;GO92(^5<E1=_/7E-5R4CD(2Z#H4-
aETAF4XKQ4Z1IVV/U.7W><H14aaBR.)](^QV,g(OI?0BY?WO4e]H+e9XTFCd5a37
b,f+cC[R3W?TY;]L/dP&3&f/A[.8HeTLRW/&FI:#1ROe<LZ)>-SW6/R&K1<eMX^]
<Z,.7[2C[Z74DgJ0IfM-?U;_02GSR5\9Y9UW<=)N+>g4f]3fM2<[T-d3(F#_P6XH
H/-bNFO)[PVRM_@L>36H.8R,fK@ge4+Y<+;H1b9O2S=>ee5;aOESdS,9,.5f?4e;
N&5[CHeK5NV3G>=6Me/;_7)TBe>G@W)#)>gR,>V5Z4&78Nd8/1?cG0VBHVWSS:6(
_:VLIQFC\-(DTE#>A4#cJf];d>VN8X7<6[D.f[f\IZ6X7YVN,3FWAGA[7eGbc:^;
D^:ZfP54,WK#TZ5A86>XU(5_[LPBY5[RK@1QP6J.)g,+YP[52\(#:_WA<A5Aa0dC
8.O0]_Q>A(c]C6O--ETC<>G9CR(AeEICAbIbOI2(\e<ZaC)fN:Q086D[R&,Q@M&Z
U,?[+0;S&<T/7Z2>XOG^R8PYW>,H;#ScDJZX2I5_=<a#Q7,KENM2J53WR?gO4D>&
Xe6FWc=DfNP<fZOd&)D<.TS\:HQ=MX)<1YV\g5VR6S<a?QHU;ACdV:9@3<M+?d+:
:1GQ=IJDU)=aYUdUWKD#&LPB]d,A>&?<K(Z/9._P&Y81fGS^M[93C;>(_gce]]G2
2XJd=WECSg@5g\4eGXCW_K=7(C6[G#IV8#+C+(WEVI;7RWN.U\SAP_R<YK:BLVI3
H^70bKLN<N8=;Wedd/bagE)3FUeB)?R8R0.ILTDU[MSS^4S.G5&JQ2R/.HABc@TH
@dQA#W<)B\b\0+H_M&Hc=(:WINbK_4(N25P6Y#RIc;ED/(LA,LdB^ERHSV<;F)L+
WIGDb_MU8SST@a>YCJ?e)XPODg;<.8L2b-7Y^?eC>,LT.0IV>(D2,W7A9R@7PZ^T
AVJbFQD?&AJL<.S7/)g\/7>5PJggOB]\EK.R^W[MJdF+)GT@ef@=)bgV:,Y&Je^[
P4d@dK,X.SAcS4+7)?^VQGd2Jc9X(MN-,V)W;a1<2dM(T8WOI>&6D93f8d&<+XIf
)+1JK8SeP_CgeD?T=9.G9\27gUXV?b@^+4=]3#cGR;N_a\fB2F2MHF8\H5G1G-4I
L]?E1FN58B.A9UL[:/@EUJ;S#9.T(,#UN-61\MRb)N^R&F^-HEB[<QTMHH)<\b:)
0+=;aAba/fGacB0f72-=F?@0ae/B9A.:X2aAPUSN75-(3;gK#d[4B;Y7?2_=^2NS
2d2UTP<.T)Z[?FbI=6E,I<HG1V9.TG\Uc?>4OFIcX\M-LIVM@514E(A,:+/\_Rg6
=-9CM6WU:ZL?B\DFXB,cO=d^+6<OS+f-OKZe==-_.YP1BN+D[Z7.S=-WQSD:WQCG
@^)]HE:?C.XOW]6Ye_B9DKME_&,#<[7V/Gb/b<-)>:LATbg<7L@YBB?+@]2N4GG;
C9EcZH?I60?XH+5bI>T@41bP0G^0N,QCd>0+_-GH\#cUEaT2P.2_(K8GR>^LX07X
<AN=K)c9)2:O/fS\_0JH0VX4[8UFbM.8YY5I&T=.b[_ULbd5EPMR\@7>=TK^cX1(
_&5g9U8M)?C(D0(:./UC4U;]5PENB>0[N?5QIR6J]YAT>+-g<\1O,S.)WVEQI[FD
LWBFRW9M^I@N>_8MU_FL&2\eA[UTKeC.4BF&fgRPV&_PaW_:gV1Q;RBc2U3#[>F[
N?QC5E3b.4]\3##3\9,E)VW?UCV2NM[aC;&9cI<(.cPc_((;Fga2[CRAH3\>XG07
V6UP2C<8&&bD^ECc21\7VC;L0b(KQ:2YOQ.S8fS+IE@0MCAc3_W>;_F?^[a&K,0>
a=f.Z1&M?b(#_,UFZI).f&(bU,3QM^./E?/QPDG/g-PD2R1N0?a;5&G>U@A)I:-,
4LCA)/6ASM-?])D8>,cc[_/5eWQdWb-;c)N&Z]3C182W(?&I#ZMV.,>AB9IgJTDQ
<13G:PU5MD.#UeMW903+P[G\+CcH>XK#K2L&WCVI2gWQ_5N]LL26D0C+1Q5&\5Wc
,:4Tb>^G41+a;91YdF@OQ33T_[2:GZ@^:;#bWb=Y#GT?,ID6fJ@Y;>A,&-XATf:5
78IK.<H043EcT193L^Wg_eP/W.8]\-L.()[Q-9JTF.7eXX?#JQ+Pfe>cOYR\LY=-
L2;#UBJ+eZ2Jc#Z0PDNMD3-3Z6Z_KN;AS9C(aIW;1<fKW=6T3&2D#(^8_\-3D90Y
#)H@V-Gg\(7W?;TSS;J7-3PP.82=YL:EKc2P@>U\YO;AP@617H>,EI^7g#@36\f&
6JR4e87IKOJG87;d:.-3,2W8C0\\Y.VeM\.^-FO;?,d]OMe?PZNE&I&(D.+2V3C=
[GIb+=,.Y\/15S]KL.30=+LGLC)#X&U=(e1X+U(EB=(fZ5#I8LJR(KWTX]8I2g^e
c7]c38d@<./T(-MD&.gI98]Tca/7@N83;.VA1I#O3F.<[ZY,3[,\IV34OV71.##F
.]Kd=&]D3[cN0BWRU+@(9K\D[;a=/6PJC4EC9cXb(3_]O8WU(B^>Q3(QP:(W\9)A
@FdLXP5?Y6HJI1/P]2WW5QE[#T<]W_DRc1g\(PB2]>Gb)9BYKB^_I3,AK=eFN,+6
:[D[D7gGG-Ue#LP+1&e)9aI?QbaNN6)_F5<8L_L4LJU_J4E>OC2^7D9g+2KG8gF:
_G7;N@Y^:XIZ6G=4.F[;#18QGZ@M,=T?bK9MZ5\L8IJ4>Z<I]Y=6HdQf2HI=a#Q4
c^GUd[bI/3)17]R<7f6&6/:TN#a2c\)5KS=KW4>,0U[UKA7S-1BLR=#@R^4B&(#7
ZP[f@=:/Q66M5>gWP0L82R&+&A8Lc9829;+,]V)O/d7GWaNFN3Y]O&-Y+[2:2/[e
BXaL+^=8C:.O_67)&440,+D9FO;U@;@HMG]X24>f/Y^Qg8B<7NBMIa68-@05A7#?
_GGC:TKOeD21\\-aOZ4^R.WRL\07UaI]3b\g_87gWV7:FGb3cI2f8??K:BYJ=a8O
Of7]Saf]B_3A/I5O>&[^ODXT/0WTT[@WUUU^cA]C<\RSFTf1[=_R+MeY5O;d\;09
55=T3P+WW8&O:W&>[b1EZ#VWAL==E6>3aL61#XO]d#<9)RPCEZg(M@eC(USG-E@9
efgTfdMSE2E0/\\^+_GKM-;#E#6>/@gW__83-CB+Id-7ZN9/M.Nb<\T=<(S3G[;J
O8_b3.^I1RgVGK<RM[.O6XQ]C5_;5D\69dIUW3?\/bCA8AYVV13&6c2E)H.-We<_
MI(cA3+W01>#X_VO\Wd_cNaGX2>@7L[Q]K2QKd2XGZ_ZE)aC_.8.BJ8Y<>,G)_9<
\?ZHBQXTKeO)cN:,C::g5A&7((3J2/W0RB@;8,dX,2_a/>e>98X[3/W0HKbD<S@+
ac6=HD-<X@WbCRHZ-UD15g41,5e;Fe2[HgdTO@,@@D_1\>2#IG9@(?c.9()YV;&]
C<;Je,XG<_R-P(VIT3;Pg((:gF]-2J_LXO.PG=gK&W8fRK1;8@9.TIU(S&BV;O<5
NA1HI+RP=2H^F)FIR\0bO)_eC[G&;G_1)P;Nf(4TP#I.RQ-R;L5G2NLE?K0;,/6f
eXJZ2cF4P@SfQXV1,Q0R7EU7&M,B6FS73H_S]C,R5-M><,8Kcd+PM=ZfB#U=R?/<
GUe)a11WIBH]aD8B)_/3@+,:f9LZJ0S>?K8g.E7g7:?,2U-Oa_9Jb+LPTd+?;QO&
,Qb_0F4M5:\]NX;:;.BBSfVf9SMM5S2FAD]G)2c7aUVEf.d4Ae;Z6abL1FM=N]<>
ObZ+0Z@#_5U1f1ZbO/<g?N[S@MU+E5G2F9.4&.V-)E;S[bBNb0Y.UY8RLQcK]SO6
Y7FJB\=2\HV9_?3S<@?^Kf84<914=<6?d.0AW;GKDGA&ff/OPGAJ^8YB+Bf-;6//
E8JH);:dNF.9SOS@3G^3cR:K5Z0+0F_\]/=.7M3R7\N;/5IM)/C\&O)B>ba7N#aF
P1Z>b-P_[H8.)^A+^(64P^7&EfMLA/3OcG2PQS2;fD/M(JEZFgPPe3213^HDXTc&
8Xf-MN=C_>=(G,?+NPcQORVI2GPNDeb6?Ba=A(BHCS?P+N)E;_,g<)dRcU^eBb/2
+a^-O7=ZML:/0-aCfLFLA-a#YL@V);]L0APSGL#68FB>_7PUV8eTWU_gQ;24K<&=
;6OQ&fce]62G#4>U\-_J6T_L?]=\gF(aW;ZQ[@9>30,6S8gE,#[Q@M-2[7Pd481g
V-dB1>GN]LK@1.N2R:M9;H@?VU2-?FaJMP/J,\;\8G)^a^3B7V:d5H_7VL/2WI4^
89T2@a3;3L,GI2\FU=[/@.T<WL7>+,]e8;U-XN.=1S=?H]F17;[9-,aGRC\JTbWS
<.>d:DJ-H^Q+Qb,d5&O-J_]?F5GdF<IJ8bGXOdKI;O<\2/&U&V?XSA]F-)cTM/@E
CR<4&L^,XQT,VaAXV2L^I_/+QRB?4#J2d_A:LU^7#X_6&\&=&_+VTSA.#ADBXZZ>
:L)_M]SPY&=Y5Z-)V-VHXQ,IHbf<+KV9)MG.,_#9ZOQEMO^CNYCcTD-bR3GQKf@=
5/bHMCH8?c@,R,3B[;;Pa+Y?MG_(LbfKL&KG)>#/BKbf8<?#c6315Afb5Ng9LCH\
1,KY(T>^Yf8<EEWF&Z/ZQFL5Z]OKN5&:S.Hcb<.RT(@0Q+^V@.4aGGfg7a)^_TYD
:ZH(_b41.L5;JH#J_D,Z6MOe&I47d9L7d[ge#cgN6gU1M;@3P<+.U)=PJPDCf3=E
1+VTS_bc+2Q(^cB1:c(E.3P=IEPGVMQ1bT2FCY;J)AV#5B2[UHMD89L\P=M3Z^T@
79dSaN2:DC?^MM5EUI:/MG_0cQG?A,OK,L(,JDD;/KbM/\_g2@AVG8R8C-+,9gI/
VL/>^93g5JASRYMLV\<1HFgB3C.3@;)>HZgPa5#cOD2]_\Z^0L>U=;gTGA1,[\bg
=@^+7eb&N<4?Y_C9-fV1B:a##W3[0f;^/-)W@OZ[]Q8M+;(86SPJ][6^(6AE\^5P
Q=<)A1DVB9>AY8G@5(>2J=R(R7;6-:EIdfP#[bDVXdQF:aAJG1GO6OCS\gNe_Y=_
<R\CCR6Gd&aROCZ[L[<<,9/DP(4-aHC99KD2:-JaNK#>J()W@[>f1Nd^R(7S6LG2
GKD<YL,&TX/B6.+G_@5IZF<b<),YRGVFL3Z]T?F(=CU@6:@#VH?;eM:W_d.63TEV
G)Q\cUag@=QH#Wa@4)AJFd1L6fU>ICO+#T7\Ea^?_PX.3e&1&F:[\IV3CYZ-CSEY
ES.H]cGXRA,(78CQI>Zd+)=b-5UI_#@NfFY)LcF^>9)T?JXK+d6+]4G@bXG7)^>J
@YTJ#_TceD6-9gYSAN(/-69S1fQg((8M@6,+3^gXQ@4NI&:f:;He8M7XDTP)Z,:<
bQLb.>,4P,.:a02\5A)./3U@4)eRI_/(;^TQP^-D2FLT_d])9+d_bAOD9KB@fSRZ
=/68H3dP?T(IEe9f)_5X@F<_X_eK=eK5)6c\D021\MT+;-f?6^Ka+Mdd2PS&DBge
)FT++J2-1#6QTUN&\-I#>6N5,cN,_M4SFZ#a?.106\b_d],=N[JPafDF^bH_HTB(
ac<?gFJ)<N>NBNK30NbSHdCbAH2,]=J=aTQb5M40A6N_8b;d/0.e;;MC&SG<;AUV
6?9C-NKX^?.e\:9[:E->50,N(09TM,HTIFZ50Vb+9C)K#79&\R7TC#)V&ILUX]YH
9B76VTHg4)XPW+]<+IZ_bZMAg<IOQdNZ9&]J+d3[,Y([2UGB:OT#GXGHMPR].]Q7
(<+.b&\9H?/cU6,1eP>O5/I&O-V2PK&J(\>/7@8\?\YLVPAULYKG\IBDZ6]bT+BH
Yd1-B1O)@-HKC/c:,D?c?M.Y2D_WQ3Zb/.1IPaB-S2EVOL.:dA3STUZKLQ&E0A\(
VEVI1PXRMg&PGUZ^I=7-)=&_+)8fYI,H4I?[:Kb00D#:)?/Q-FFYAO^cg/LS4TLG
E7J=E=MDXPR2H4QBA,]g5aI8UZdc>f(TEG_TB/aES-NJ@\e+_5T/H_beVQ]L-d#^
ZOBd3J_<K=[HX#D,?0G/EL[_g.BMKX7R\f(7MUY>5=X#eBFW3DafHNL[;8S,1K^&
S-H9BHHGIG4@[a(8f&3@R964JHMC5YHM=0)_HHS]07GD^^):8/@C2AN:C3[/9Uc:
514EB2B9XB4,b6[GM@\9J1(cSK]D./E-]MG:JPRd:_K_=d.Sd.EfB4@:+caP?c<@
=>ZJ76d1b2#+acE.&#>We[.A,&;BECaO<L+g[;8_gR<L@(Ae5#<&ebgM?AZ3R-Y4
P,_(+C5-B#/FMQTd9M=8cI;3L_3NWB?Be^Jge(IC6O9^[>]\TTOTCdSPALYIaYK)
I-80-.X+)3(;dR7PW@BUCCc.MZcLg;>F&Nd8W1H#NgLAALOT:\#dL;IgX6)#PN[&
dJ,)be&bLAN#ED6=VDKJ)-G89/1M<LE&K)c?2AgSN8+O&T-=fRC[^?&E,#,?+.PV
&Q_Z(dI8V7cTZ4J_3RG8&N>@)R9,^7J?BMHK-\M2[O9M\)03Z1W@>L;+ETSF;<a/
+43NR)NMb>R:>4JB8Ub9&4/KM1-<<2]9DGSBgeAa?-V0WJ-4.]1Ic\-Y2K@F]YB-
AS(Jd(9cM_X.eIZANbKc]^GP6U^J5eI_ZY_-bXX)7SAZU\NT>VV@fXCZWV?N:IW&
_dReTF^883QJgV#2.P@)KFaa,g?EP=HBa\&:A+,N_.K3K4696CC=GD4N8_f]7a_X
OAgP9(b\[?_g,T9;Af[e[D724^PTA#I.fa<WIS2+Sa6Z&=JYBPAA5HX+1JE<(\gH
M9/5^8.D?MPf&_7bde8M@DAdK/J>R;MGBW3[4.:1IC_/\R3?]a8#3/5+]4CZ1cD)
BWN34M1+6B]NZ<]_A550(2S(3eN23-6E27M.?X-C&ReD&_e(3:M^WbXU8[bVAU5E
<_IM7G;bP_.\OBA(04D&98^b&e5NIB6dAWGde0E:b/aGJ)G1U<SZ@Bb,gSXNMTC:
7J@K<[XAM]NX0IbRQXgEd;_:O5b4Ggd.2\?R:DCd/QB8:5eTDH6\T1NLUE(,N1<J
c-E@,&<&G@<3WXO&DSB,^?/3/a\3<E2(;T1Mb^&FLWQA/d(#]3<?G)@2PVc;c6/O
2]T,9O?#CGT;;+9?K<S>[,?2-SK;bK4UE/N+TFTOe\APS:YABA8-6V8VE#]dQ5dd
UWW[;eLSK4Q&WD,cUS9Vf[QKIgWd(,e^=?B_Ub08-/bXEKT)c?d=.d/_\CHD[;c9
-dUb=ML;6M>gN??>F<BC7Q@05P18P.N;S[9A<QAQaXMM3GQC-g:8cM&cGA<DM5:L
:+X]_@QcB7f+NeQQ\E/TdC&X&41:@PT:#]SH4:IJ[[8#E<Y[O20=+E5g2):,_894
C@;TCI,H4D/<S+0VA<GV7WQ^J@6,#A->.X?Q6eMD[a4P72/e#.=Yc]A<VLTT(Ef,
KPcHS916&UY6XA>:X=HgGC?b-bd@[<9.IG<NJ^(eA\_@[NQ_aF3]JIfB>HZ2<f/^
R&+8#-C>DbUF4=OQ22X3)gC[:RC[7+[Q#:,PI2]SR&H+>-UJ#]VO4>NU3Q<JGB^:
73Q7=A8LO1b4dZ5[8+?#b)f0-?53MU(8A+cbN:gB@,)c/4-RQ-]bZ:K=eM(I#f<e
#Y7X5-B6CJ34,$
`endprotected
endmodule